library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
library unisim;
use unisim.vcomponents.all;

--############################################################################--
--#                       File generated automatically                       #--
--#                            by inst_muxes.py                              #--
--#                                                                          #--
--#                python inst_muxes.py > mii_shifter_lut.vhd                #--
--############################################################################--


entity mii_shifter_lut is
  Port(
    in_0      : in std_logic_vector(255 downto 0);
    in_1      : in std_logic_vector(255 downto 0);
    sel_mux   : in std_logic_vector(2 downto 0);

    data_out  : out std_logic_vector(255 downto 0)
  );
end entity;


architecture behav_mii_shifter of mii_shifter_lut is
  component mux8 is
    Port (  data_in : in std_logic_vector(7 downto 0);
                sel : in std_logic_vector(2 downto 0);
           data_out : out std_logic
          );
  end component;
-- Signal declarations:
signal mux_input_0 : std_logic_vector(7 downto 0);
signal mux_input_1 : std_logic_vector(7 downto 0);
signal mux_input_2 : std_logic_vector(7 downto 0);
signal mux_input_3 : std_logic_vector(7 downto 0);
signal mux_input_4 : std_logic_vector(7 downto 0);
signal mux_input_5 : std_logic_vector(7 downto 0);
signal mux_input_6 : std_logic_vector(7 downto 0);
signal mux_input_7 : std_logic_vector(7 downto 0);
signal mux_input_8 : std_logic_vector(7 downto 0);
signal mux_input_9 : std_logic_vector(7 downto 0);
signal mux_input_10 : std_logic_vector(7 downto 0);
signal mux_input_11 : std_logic_vector(7 downto 0);
signal mux_input_12 : std_logic_vector(7 downto 0);
signal mux_input_13 : std_logic_vector(7 downto 0);
signal mux_input_14 : std_logic_vector(7 downto 0);
signal mux_input_15 : std_logic_vector(7 downto 0);
signal mux_input_16 : std_logic_vector(7 downto 0);
signal mux_input_17 : std_logic_vector(7 downto 0);
signal mux_input_18 : std_logic_vector(7 downto 0);
signal mux_input_19 : std_logic_vector(7 downto 0);
signal mux_input_20 : std_logic_vector(7 downto 0);
signal mux_input_21 : std_logic_vector(7 downto 0);
signal mux_input_22 : std_logic_vector(7 downto 0);
signal mux_input_23 : std_logic_vector(7 downto 0);
signal mux_input_24 : std_logic_vector(7 downto 0);
signal mux_input_25 : std_logic_vector(7 downto 0);
signal mux_input_26 : std_logic_vector(7 downto 0);
signal mux_input_27 : std_logic_vector(7 downto 0);
signal mux_input_28 : std_logic_vector(7 downto 0);
signal mux_input_29 : std_logic_vector(7 downto 0);
signal mux_input_30 : std_logic_vector(7 downto 0);
signal mux_input_31 : std_logic_vector(7 downto 0);
signal mux_input_32 : std_logic_vector(7 downto 0);
signal mux_input_33 : std_logic_vector(7 downto 0);
signal mux_input_34 : std_logic_vector(7 downto 0);
signal mux_input_35 : std_logic_vector(7 downto 0);
signal mux_input_36 : std_logic_vector(7 downto 0);
signal mux_input_37 : std_logic_vector(7 downto 0);
signal mux_input_38 : std_logic_vector(7 downto 0);
signal mux_input_39 : std_logic_vector(7 downto 0);
signal mux_input_40 : std_logic_vector(7 downto 0);
signal mux_input_41 : std_logic_vector(7 downto 0);
signal mux_input_42 : std_logic_vector(7 downto 0);
signal mux_input_43 : std_logic_vector(7 downto 0);
signal mux_input_44 : std_logic_vector(7 downto 0);
signal mux_input_45 : std_logic_vector(7 downto 0);
signal mux_input_46 : std_logic_vector(7 downto 0);
signal mux_input_47 : std_logic_vector(7 downto 0);
signal mux_input_48 : std_logic_vector(7 downto 0);
signal mux_input_49 : std_logic_vector(7 downto 0);
signal mux_input_50 : std_logic_vector(7 downto 0);
signal mux_input_51 : std_logic_vector(7 downto 0);
signal mux_input_52 : std_logic_vector(7 downto 0);
signal mux_input_53 : std_logic_vector(7 downto 0);
signal mux_input_54 : std_logic_vector(7 downto 0);
signal mux_input_55 : std_logic_vector(7 downto 0);
signal mux_input_56 : std_logic_vector(7 downto 0);
signal mux_input_57 : std_logic_vector(7 downto 0);
signal mux_input_58 : std_logic_vector(7 downto 0);
signal mux_input_59 : std_logic_vector(7 downto 0);
signal mux_input_60 : std_logic_vector(7 downto 0);
signal mux_input_61 : std_logic_vector(7 downto 0);
signal mux_input_62 : std_logic_vector(7 downto 0);
signal mux_input_63 : std_logic_vector(7 downto 0);
signal mux_input_64 : std_logic_vector(7 downto 0);
signal mux_input_65 : std_logic_vector(7 downto 0);
signal mux_input_66 : std_logic_vector(7 downto 0);
signal mux_input_67 : std_logic_vector(7 downto 0);
signal mux_input_68 : std_logic_vector(7 downto 0);
signal mux_input_69 : std_logic_vector(7 downto 0);
signal mux_input_70 : std_logic_vector(7 downto 0);
signal mux_input_71 : std_logic_vector(7 downto 0);
signal mux_input_72 : std_logic_vector(7 downto 0);
signal mux_input_73 : std_logic_vector(7 downto 0);
signal mux_input_74 : std_logic_vector(7 downto 0);
signal mux_input_75 : std_logic_vector(7 downto 0);
signal mux_input_76 : std_logic_vector(7 downto 0);
signal mux_input_77 : std_logic_vector(7 downto 0);
signal mux_input_78 : std_logic_vector(7 downto 0);
signal mux_input_79 : std_logic_vector(7 downto 0);
signal mux_input_80 : std_logic_vector(7 downto 0);
signal mux_input_81 : std_logic_vector(7 downto 0);
signal mux_input_82 : std_logic_vector(7 downto 0);
signal mux_input_83 : std_logic_vector(7 downto 0);
signal mux_input_84 : std_logic_vector(7 downto 0);
signal mux_input_85 : std_logic_vector(7 downto 0);
signal mux_input_86 : std_logic_vector(7 downto 0);
signal mux_input_87 : std_logic_vector(7 downto 0);
signal mux_input_88 : std_logic_vector(7 downto 0);
signal mux_input_89 : std_logic_vector(7 downto 0);
signal mux_input_90 : std_logic_vector(7 downto 0);
signal mux_input_91 : std_logic_vector(7 downto 0);
signal mux_input_92 : std_logic_vector(7 downto 0);
signal mux_input_93 : std_logic_vector(7 downto 0);
signal mux_input_94 : std_logic_vector(7 downto 0);
signal mux_input_95 : std_logic_vector(7 downto 0);
signal mux_input_96 : std_logic_vector(7 downto 0);
signal mux_input_97 : std_logic_vector(7 downto 0);
signal mux_input_98 : std_logic_vector(7 downto 0);
signal mux_input_99 : std_logic_vector(7 downto 0);
signal mux_input_100 : std_logic_vector(7 downto 0);
signal mux_input_101 : std_logic_vector(7 downto 0);
signal mux_input_102 : std_logic_vector(7 downto 0);
signal mux_input_103 : std_logic_vector(7 downto 0);
signal mux_input_104 : std_logic_vector(7 downto 0);
signal mux_input_105 : std_logic_vector(7 downto 0);
signal mux_input_106 : std_logic_vector(7 downto 0);
signal mux_input_107 : std_logic_vector(7 downto 0);
signal mux_input_108 : std_logic_vector(7 downto 0);
signal mux_input_109 : std_logic_vector(7 downto 0);
signal mux_input_110 : std_logic_vector(7 downto 0);
signal mux_input_111 : std_logic_vector(7 downto 0);
signal mux_input_112 : std_logic_vector(7 downto 0);
signal mux_input_113 : std_logic_vector(7 downto 0);
signal mux_input_114 : std_logic_vector(7 downto 0);
signal mux_input_115 : std_logic_vector(7 downto 0);
signal mux_input_116 : std_logic_vector(7 downto 0);
signal mux_input_117 : std_logic_vector(7 downto 0);
signal mux_input_118 : std_logic_vector(7 downto 0);
signal mux_input_119 : std_logic_vector(7 downto 0);
signal mux_input_120 : std_logic_vector(7 downto 0);
signal mux_input_121 : std_logic_vector(7 downto 0);
signal mux_input_122 : std_logic_vector(7 downto 0);
signal mux_input_123 : std_logic_vector(7 downto 0);
signal mux_input_124 : std_logic_vector(7 downto 0);
signal mux_input_125 : std_logic_vector(7 downto 0);
signal mux_input_126 : std_logic_vector(7 downto 0);
signal mux_input_127 : std_logic_vector(7 downto 0);
signal mux_input_128 : std_logic_vector(7 downto 0);
signal mux_input_129 : std_logic_vector(7 downto 0);
signal mux_input_130 : std_logic_vector(7 downto 0);
signal mux_input_131 : std_logic_vector(7 downto 0);
signal mux_input_132 : std_logic_vector(7 downto 0);
signal mux_input_133 : std_logic_vector(7 downto 0);
signal mux_input_134 : std_logic_vector(7 downto 0);
signal mux_input_135 : std_logic_vector(7 downto 0);
signal mux_input_136 : std_logic_vector(7 downto 0);
signal mux_input_137 : std_logic_vector(7 downto 0);
signal mux_input_138 : std_logic_vector(7 downto 0);
signal mux_input_139 : std_logic_vector(7 downto 0);
signal mux_input_140 : std_logic_vector(7 downto 0);
signal mux_input_141 : std_logic_vector(7 downto 0);
signal mux_input_142 : std_logic_vector(7 downto 0);
signal mux_input_143 : std_logic_vector(7 downto 0);
signal mux_input_144 : std_logic_vector(7 downto 0);
signal mux_input_145 : std_logic_vector(7 downto 0);
signal mux_input_146 : std_logic_vector(7 downto 0);
signal mux_input_147 : std_logic_vector(7 downto 0);
signal mux_input_148 : std_logic_vector(7 downto 0);
signal mux_input_149 : std_logic_vector(7 downto 0);
signal mux_input_150 : std_logic_vector(7 downto 0);
signal mux_input_151 : std_logic_vector(7 downto 0);
signal mux_input_152 : std_logic_vector(7 downto 0);
signal mux_input_153 : std_logic_vector(7 downto 0);
signal mux_input_154 : std_logic_vector(7 downto 0);
signal mux_input_155 : std_logic_vector(7 downto 0);
signal mux_input_156 : std_logic_vector(7 downto 0);
signal mux_input_157 : std_logic_vector(7 downto 0);
signal mux_input_158 : std_logic_vector(7 downto 0);
signal mux_input_159 : std_logic_vector(7 downto 0);
signal mux_input_160 : std_logic_vector(7 downto 0);
signal mux_input_161 : std_logic_vector(7 downto 0);
signal mux_input_162 : std_logic_vector(7 downto 0);
signal mux_input_163 : std_logic_vector(7 downto 0);
signal mux_input_164 : std_logic_vector(7 downto 0);
signal mux_input_165 : std_logic_vector(7 downto 0);
signal mux_input_166 : std_logic_vector(7 downto 0);
signal mux_input_167 : std_logic_vector(7 downto 0);
signal mux_input_168 : std_logic_vector(7 downto 0);
signal mux_input_169 : std_logic_vector(7 downto 0);
signal mux_input_170 : std_logic_vector(7 downto 0);
signal mux_input_171 : std_logic_vector(7 downto 0);
signal mux_input_172 : std_logic_vector(7 downto 0);
signal mux_input_173 : std_logic_vector(7 downto 0);
signal mux_input_174 : std_logic_vector(7 downto 0);
signal mux_input_175 : std_logic_vector(7 downto 0);
signal mux_input_176 : std_logic_vector(7 downto 0);
signal mux_input_177 : std_logic_vector(7 downto 0);
signal mux_input_178 : std_logic_vector(7 downto 0);
signal mux_input_179 : std_logic_vector(7 downto 0);
signal mux_input_180 : std_logic_vector(7 downto 0);
signal mux_input_181 : std_logic_vector(7 downto 0);
signal mux_input_182 : std_logic_vector(7 downto 0);
signal mux_input_183 : std_logic_vector(7 downto 0);
signal mux_input_184 : std_logic_vector(7 downto 0);
signal mux_input_185 : std_logic_vector(7 downto 0);
signal mux_input_186 : std_logic_vector(7 downto 0);
signal mux_input_187 : std_logic_vector(7 downto 0);
signal mux_input_188 : std_logic_vector(7 downto 0);
signal mux_input_189 : std_logic_vector(7 downto 0);
signal mux_input_190 : std_logic_vector(7 downto 0);
signal mux_input_191 : std_logic_vector(7 downto 0);
signal mux_input_192 : std_logic_vector(7 downto 0);
signal mux_input_193 : std_logic_vector(7 downto 0);
signal mux_input_194 : std_logic_vector(7 downto 0);
signal mux_input_195 : std_logic_vector(7 downto 0);
signal mux_input_196 : std_logic_vector(7 downto 0);
signal mux_input_197 : std_logic_vector(7 downto 0);
signal mux_input_198 : std_logic_vector(7 downto 0);
signal mux_input_199 : std_logic_vector(7 downto 0);
signal mux_input_200 : std_logic_vector(7 downto 0);
signal mux_input_201 : std_logic_vector(7 downto 0);
signal mux_input_202 : std_logic_vector(7 downto 0);
signal mux_input_203 : std_logic_vector(7 downto 0);
signal mux_input_204 : std_logic_vector(7 downto 0);
signal mux_input_205 : std_logic_vector(7 downto 0);
signal mux_input_206 : std_logic_vector(7 downto 0);
signal mux_input_207 : std_logic_vector(7 downto 0);
signal mux_input_208 : std_logic_vector(7 downto 0);
signal mux_input_209 : std_logic_vector(7 downto 0);
signal mux_input_210 : std_logic_vector(7 downto 0);
signal mux_input_211 : std_logic_vector(7 downto 0);
signal mux_input_212 : std_logic_vector(7 downto 0);
signal mux_input_213 : std_logic_vector(7 downto 0);
signal mux_input_214 : std_logic_vector(7 downto 0);
signal mux_input_215 : std_logic_vector(7 downto 0);
signal mux_input_216 : std_logic_vector(7 downto 0);
signal mux_input_217 : std_logic_vector(7 downto 0);
signal mux_input_218 : std_logic_vector(7 downto 0);
signal mux_input_219 : std_logic_vector(7 downto 0);
signal mux_input_220 : std_logic_vector(7 downto 0);
signal mux_input_221 : std_logic_vector(7 downto 0);
signal mux_input_222 : std_logic_vector(7 downto 0);
signal mux_input_223 : std_logic_vector(7 downto 0);
signal mux_input_224 : std_logic_vector(7 downto 0);
signal mux_input_225 : std_logic_vector(7 downto 0);
signal mux_input_226 : std_logic_vector(7 downto 0);
signal mux_input_227 : std_logic_vector(7 downto 0);
signal mux_input_228 : std_logic_vector(7 downto 0);
signal mux_input_229 : std_logic_vector(7 downto 0);
signal mux_input_230 : std_logic_vector(7 downto 0);
signal mux_input_231 : std_logic_vector(7 downto 0);
signal mux_input_232 : std_logic_vector(7 downto 0);
signal mux_input_233 : std_logic_vector(7 downto 0);
signal mux_input_234 : std_logic_vector(7 downto 0);
signal mux_input_235 : std_logic_vector(7 downto 0);
signal mux_input_236 : std_logic_vector(7 downto 0);
signal mux_input_237 : std_logic_vector(7 downto 0);
signal mux_input_238 : std_logic_vector(7 downto 0);
signal mux_input_239 : std_logic_vector(7 downto 0);
signal mux_input_240 : std_logic_vector(7 downto 0);
signal mux_input_241 : std_logic_vector(7 downto 0);
signal mux_input_242 : std_logic_vector(7 downto 0);
signal mux_input_243 : std_logic_vector(7 downto 0);
signal mux_input_244 : std_logic_vector(7 downto 0);
signal mux_input_245 : std_logic_vector(7 downto 0);
signal mux_input_246 : std_logic_vector(7 downto 0);
signal mux_input_247 : std_logic_vector(7 downto 0);
signal mux_input_248 : std_logic_vector(7 downto 0);
signal mux_input_249 : std_logic_vector(7 downto 0);
signal mux_input_250 : std_logic_vector(7 downto 0);
signal mux_input_251 : std_logic_vector(7 downto 0);
signal mux_input_252 : std_logic_vector(7 downto 0);
signal mux_input_253 : std_logic_vector(7 downto 0);
signal mux_input_254 : std_logic_vector(7 downto 0);
signal mux_input_255 : std_logic_vector(7 downto 0);
begin
-- Muxes from 0 to 31:
mux_input_0 <= in_1(224) & in_1(192) & in_1(160) & in_1(128) & in_1(96) & in_1(64) & in_1(32) & in_1(0);
mux_input_1 <= in_1(225) & in_1(193) & in_1(161) & in_1(129) & in_1(97) & in_1(65) & in_1(33) & in_1(1);
mux_input_2 <= in_1(226) & in_1(194) & in_1(162) & in_1(130) & in_1(98) & in_1(66) & in_1(34) & in_1(2);
mux_input_3 <= in_1(227) & in_1(195) & in_1(163) & in_1(131) & in_1(99) & in_1(67) & in_1(35) & in_1(3);
mux_input_4 <= in_1(228) & in_1(196) & in_1(164) & in_1(132) & in_1(100) & in_1(68) & in_1(36) & in_1(4);
mux_input_5 <= in_1(229) & in_1(197) & in_1(165) & in_1(133) & in_1(101) & in_1(69) & in_1(37) & in_1(5);
mux_input_6 <= in_1(230) & in_1(198) & in_1(166) & in_1(134) & in_1(102) & in_1(70) & in_1(38) & in_1(6);
mux_input_7 <= in_1(231) & in_1(199) & in_1(167) & in_1(135) & in_1(103) & in_1(71) & in_1(39) & in_1(7);
mux_input_8 <= in_1(232) & in_1(200) & in_1(168) & in_1(136) & in_1(104) & in_1(72) & in_1(40) & in_1(8);
mux_input_9 <= in_1(233) & in_1(201) & in_1(169) & in_1(137) & in_1(105) & in_1(73) & in_1(41) & in_1(9);
mux_input_10 <= in_1(234) & in_1(202) & in_1(170) & in_1(138) & in_1(106) & in_1(74) & in_1(42) & in_1(10);
mux_input_11 <= in_1(235) & in_1(203) & in_1(171) & in_1(139) & in_1(107) & in_1(75) & in_1(43) & in_1(11);
mux_input_12 <= in_1(236) & in_1(204) & in_1(172) & in_1(140) & in_1(108) & in_1(76) & in_1(44) & in_1(12);
mux_input_13 <= in_1(237) & in_1(205) & in_1(173) & in_1(141) & in_1(109) & in_1(77) & in_1(45) & in_1(13);
mux_input_14 <= in_1(238) & in_1(206) & in_1(174) & in_1(142) & in_1(110) & in_1(78) & in_1(46) & in_1(14);
mux_input_15 <= in_1(239) & in_1(207) & in_1(175) & in_1(143) & in_1(111) & in_1(79) & in_1(47) & in_1(15);
mux_input_16 <= in_1(240) & in_1(208) & in_1(176) & in_1(144) & in_1(112) & in_1(80) & in_1(48) & in_1(16);
mux_input_17 <= in_1(241) & in_1(209) & in_1(177) & in_1(145) & in_1(113) & in_1(81) & in_1(49) & in_1(17);
mux_input_18 <= in_1(242) & in_1(210) & in_1(178) & in_1(146) & in_1(114) & in_1(82) & in_1(50) & in_1(18);
mux_input_19 <= in_1(243) & in_1(211) & in_1(179) & in_1(147) & in_1(115) & in_1(83) & in_1(51) & in_1(19);
mux_input_20 <= in_1(244) & in_1(212) & in_1(180) & in_1(148) & in_1(116) & in_1(84) & in_1(52) & in_1(20);
mux_input_21 <= in_1(245) & in_1(213) & in_1(181) & in_1(149) & in_1(117) & in_1(85) & in_1(53) & in_1(21);
mux_input_22 <= in_1(246) & in_1(214) & in_1(182) & in_1(150) & in_1(118) & in_1(86) & in_1(54) & in_1(22);
mux_input_23 <= in_1(247) & in_1(215) & in_1(183) & in_1(151) & in_1(119) & in_1(87) & in_1(55) & in_1(23);
mux_input_24 <= in_1(248) & in_1(216) & in_1(184) & in_1(152) & in_1(120) & in_1(88) & in_1(56) & in_1(24);
mux_input_25 <= in_1(249) & in_1(217) & in_1(185) & in_1(153) & in_1(121) & in_1(89) & in_1(57) & in_1(25);
mux_input_26 <= in_1(250) & in_1(218) & in_1(186) & in_1(154) & in_1(122) & in_1(90) & in_1(58) & in_1(26);
mux_input_27 <= in_1(251) & in_1(219) & in_1(187) & in_1(155) & in_1(123) & in_1(91) & in_1(59) & in_1(27);
mux_input_28 <= in_1(252) & in_1(220) & in_1(188) & in_1(156) & in_1(124) & in_1(92) & in_1(60) & in_1(28);
mux_input_29 <= in_1(253) & in_1(221) & in_1(189) & in_1(157) & in_1(125) & in_1(93) & in_1(61) & in_1(29);
mux_input_30 <= in_1(254) & in_1(222) & in_1(190) & in_1(158) & in_1(126) & in_1(94) & in_1(62) & in_1(30);
mux_input_31 <= in_1(255) & in_1(223) & in_1(191) & in_1(159) & in_1(127) & in_1(95) & in_1(63) & in_1(31);
-- Muxes from 32 to 63:
mux_input_32 <= in_0(0) & in_1(224) & in_1(192) & in_1(160) & in_1(128) & in_1(96) & in_1(64) & in_1(32);
mux_input_33 <= in_0(1) & in_1(225) & in_1(193) & in_1(161) & in_1(129) & in_1(97) & in_1(65) & in_1(33);
mux_input_34 <= in_0(2) & in_1(226) & in_1(194) & in_1(162) & in_1(130) & in_1(98) & in_1(66) & in_1(34);
mux_input_35 <= in_0(3) & in_1(227) & in_1(195) & in_1(163) & in_1(131) & in_1(99) & in_1(67) & in_1(35);
mux_input_36 <= in_0(4) & in_1(228) & in_1(196) & in_1(164) & in_1(132) & in_1(100) & in_1(68) & in_1(36);
mux_input_37 <= in_0(5) & in_1(229) & in_1(197) & in_1(165) & in_1(133) & in_1(101) & in_1(69) & in_1(37);
mux_input_38 <= in_0(6) & in_1(230) & in_1(198) & in_1(166) & in_1(134) & in_1(102) & in_1(70) & in_1(38);
mux_input_39 <= in_0(7) & in_1(231) & in_1(199) & in_1(167) & in_1(135) & in_1(103) & in_1(71) & in_1(39);
mux_input_40 <= in_0(8) & in_1(232) & in_1(200) & in_1(168) & in_1(136) & in_1(104) & in_1(72) & in_1(40);
mux_input_41 <= in_0(9) & in_1(233) & in_1(201) & in_1(169) & in_1(137) & in_1(105) & in_1(73) & in_1(41);
mux_input_42 <= in_0(10) & in_1(234) & in_1(202) & in_1(170) & in_1(138) & in_1(106) & in_1(74) & in_1(42);
mux_input_43 <= in_0(11) & in_1(235) & in_1(203) & in_1(171) & in_1(139) & in_1(107) & in_1(75) & in_1(43);
mux_input_44 <= in_0(12) & in_1(236) & in_1(204) & in_1(172) & in_1(140) & in_1(108) & in_1(76) & in_1(44);
mux_input_45 <= in_0(13) & in_1(237) & in_1(205) & in_1(173) & in_1(141) & in_1(109) & in_1(77) & in_1(45);
mux_input_46 <= in_0(14) & in_1(238) & in_1(206) & in_1(174) & in_1(142) & in_1(110) & in_1(78) & in_1(46);
mux_input_47 <= in_0(15) & in_1(239) & in_1(207) & in_1(175) & in_1(143) & in_1(111) & in_1(79) & in_1(47);
mux_input_48 <= in_0(16) & in_1(240) & in_1(208) & in_1(176) & in_1(144) & in_1(112) & in_1(80) & in_1(48);
mux_input_49 <= in_0(17) & in_1(241) & in_1(209) & in_1(177) & in_1(145) & in_1(113) & in_1(81) & in_1(49);
mux_input_50 <= in_0(18) & in_1(242) & in_1(210) & in_1(178) & in_1(146) & in_1(114) & in_1(82) & in_1(50);
mux_input_51 <= in_0(19) & in_1(243) & in_1(211) & in_1(179) & in_1(147) & in_1(115) & in_1(83) & in_1(51);
mux_input_52 <= in_0(20) & in_1(244) & in_1(212) & in_1(180) & in_1(148) & in_1(116) & in_1(84) & in_1(52);
mux_input_53 <= in_0(21) & in_1(245) & in_1(213) & in_1(181) & in_1(149) & in_1(117) & in_1(85) & in_1(53);
mux_input_54 <= in_0(22) & in_1(246) & in_1(214) & in_1(182) & in_1(150) & in_1(118) & in_1(86) & in_1(54);
mux_input_55 <= in_0(23) & in_1(247) & in_1(215) & in_1(183) & in_1(151) & in_1(119) & in_1(87) & in_1(55);
mux_input_56 <= in_0(24) & in_1(248) & in_1(216) & in_1(184) & in_1(152) & in_1(120) & in_1(88) & in_1(56);
mux_input_57 <= in_0(25) & in_1(249) & in_1(217) & in_1(185) & in_1(153) & in_1(121) & in_1(89) & in_1(57);
mux_input_58 <= in_0(26) & in_1(250) & in_1(218) & in_1(186) & in_1(154) & in_1(122) & in_1(90) & in_1(58);
mux_input_59 <= in_0(27) & in_1(251) & in_1(219) & in_1(187) & in_1(155) & in_1(123) & in_1(91) & in_1(59);
mux_input_60 <= in_0(28) & in_1(252) & in_1(220) & in_1(188) & in_1(156) & in_1(124) & in_1(92) & in_1(60);
mux_input_61 <= in_0(29) & in_1(253) & in_1(221) & in_1(189) & in_1(157) & in_1(125) & in_1(93) & in_1(61);
mux_input_62 <= in_0(30) & in_1(254) & in_1(222) & in_1(190) & in_1(158) & in_1(126) & in_1(94) & in_1(62);
mux_input_63 <= in_0(31) & in_1(255) & in_1(223) & in_1(191) & in_1(159) & in_1(127) & in_1(95) & in_1(63);
-- Muxes from 64 to 95:
mux_input_64 <= in_0(32) & in_0(0) & in_1(224) & in_1(192) & in_1(160) & in_1(128) & in_1(96) & in_1(64);
mux_input_65 <= in_0(33) & in_0(1) & in_1(225) & in_1(193) & in_1(161) & in_1(129) & in_1(97) & in_1(65);
mux_input_66 <= in_0(34) & in_0(2) & in_1(226) & in_1(194) & in_1(162) & in_1(130) & in_1(98) & in_1(66);
mux_input_67 <= in_0(35) & in_0(3) & in_1(227) & in_1(195) & in_1(163) & in_1(131) & in_1(99) & in_1(67);
mux_input_68 <= in_0(36) & in_0(4) & in_1(228) & in_1(196) & in_1(164) & in_1(132) & in_1(100) & in_1(68);
mux_input_69 <= in_0(37) & in_0(5) & in_1(229) & in_1(197) & in_1(165) & in_1(133) & in_1(101) & in_1(69);
mux_input_70 <= in_0(38) & in_0(6) & in_1(230) & in_1(198) & in_1(166) & in_1(134) & in_1(102) & in_1(70);
mux_input_71 <= in_0(39) & in_0(7) & in_1(231) & in_1(199) & in_1(167) & in_1(135) & in_1(103) & in_1(71);
mux_input_72 <= in_0(40) & in_0(8) & in_1(232) & in_1(200) & in_1(168) & in_1(136) & in_1(104) & in_1(72);
mux_input_73 <= in_0(41) & in_0(9) & in_1(233) & in_1(201) & in_1(169) & in_1(137) & in_1(105) & in_1(73);
mux_input_74 <= in_0(42) & in_0(10) & in_1(234) & in_1(202) & in_1(170) & in_1(138) & in_1(106) & in_1(74);
mux_input_75 <= in_0(43) & in_0(11) & in_1(235) & in_1(203) & in_1(171) & in_1(139) & in_1(107) & in_1(75);
mux_input_76 <= in_0(44) & in_0(12) & in_1(236) & in_1(204) & in_1(172) & in_1(140) & in_1(108) & in_1(76);
mux_input_77 <= in_0(45) & in_0(13) & in_1(237) & in_1(205) & in_1(173) & in_1(141) & in_1(109) & in_1(77);
mux_input_78 <= in_0(46) & in_0(14) & in_1(238) & in_1(206) & in_1(174) & in_1(142) & in_1(110) & in_1(78);
mux_input_79 <= in_0(47) & in_0(15) & in_1(239) & in_1(207) & in_1(175) & in_1(143) & in_1(111) & in_1(79);
mux_input_80 <= in_0(48) & in_0(16) & in_1(240) & in_1(208) & in_1(176) & in_1(144) & in_1(112) & in_1(80);
mux_input_81 <= in_0(49) & in_0(17) & in_1(241) & in_1(209) & in_1(177) & in_1(145) & in_1(113) & in_1(81);
mux_input_82 <= in_0(50) & in_0(18) & in_1(242) & in_1(210) & in_1(178) & in_1(146) & in_1(114) & in_1(82);
mux_input_83 <= in_0(51) & in_0(19) & in_1(243) & in_1(211) & in_1(179) & in_1(147) & in_1(115) & in_1(83);
mux_input_84 <= in_0(52) & in_0(20) & in_1(244) & in_1(212) & in_1(180) & in_1(148) & in_1(116) & in_1(84);
mux_input_85 <= in_0(53) & in_0(21) & in_1(245) & in_1(213) & in_1(181) & in_1(149) & in_1(117) & in_1(85);
mux_input_86 <= in_0(54) & in_0(22) & in_1(246) & in_1(214) & in_1(182) & in_1(150) & in_1(118) & in_1(86);
mux_input_87 <= in_0(55) & in_0(23) & in_1(247) & in_1(215) & in_1(183) & in_1(151) & in_1(119) & in_1(87);
mux_input_88 <= in_0(56) & in_0(24) & in_1(248) & in_1(216) & in_1(184) & in_1(152) & in_1(120) & in_1(88);
mux_input_89 <= in_0(57) & in_0(25) & in_1(249) & in_1(217) & in_1(185) & in_1(153) & in_1(121) & in_1(89);
mux_input_90 <= in_0(58) & in_0(26) & in_1(250) & in_1(218) & in_1(186) & in_1(154) & in_1(122) & in_1(90);
mux_input_91 <= in_0(59) & in_0(27) & in_1(251) & in_1(219) & in_1(187) & in_1(155) & in_1(123) & in_1(91);
mux_input_92 <= in_0(60) & in_0(28) & in_1(252) & in_1(220) & in_1(188) & in_1(156) & in_1(124) & in_1(92);
mux_input_93 <= in_0(61) & in_0(29) & in_1(253) & in_1(221) & in_1(189) & in_1(157) & in_1(125) & in_1(93);
mux_input_94 <= in_0(62) & in_0(30) & in_1(254) & in_1(222) & in_1(190) & in_1(158) & in_1(126) & in_1(94);
mux_input_95 <= in_0(63) & in_0(31) & in_1(255) & in_1(223) & in_1(191) & in_1(159) & in_1(127) & in_1(95);
-- Muxes from 96 to 127:
mux_input_96 <= in_0(64) & in_0(32) & in_0(0) & in_1(224) & in_1(192) & in_1(160) & in_1(128) & in_1(96);
mux_input_97 <= in_0(65) & in_0(33) & in_0(1) & in_1(225) & in_1(193) & in_1(161) & in_1(129) & in_1(97);
mux_input_98 <= in_0(66) & in_0(34) & in_0(2) & in_1(226) & in_1(194) & in_1(162) & in_1(130) & in_1(98);
mux_input_99 <= in_0(67) & in_0(35) & in_0(3) & in_1(227) & in_1(195) & in_1(163) & in_1(131) & in_1(99);
mux_input_100 <= in_0(68) & in_0(36) & in_0(4) & in_1(228) & in_1(196) & in_1(164) & in_1(132) & in_1(100);
mux_input_101 <= in_0(69) & in_0(37) & in_0(5) & in_1(229) & in_1(197) & in_1(165) & in_1(133) & in_1(101);
mux_input_102 <= in_0(70) & in_0(38) & in_0(6) & in_1(230) & in_1(198) & in_1(166) & in_1(134) & in_1(102);
mux_input_103 <= in_0(71) & in_0(39) & in_0(7) & in_1(231) & in_1(199) & in_1(167) & in_1(135) & in_1(103);
mux_input_104 <= in_0(72) & in_0(40) & in_0(8) & in_1(232) & in_1(200) & in_1(168) & in_1(136) & in_1(104);
mux_input_105 <= in_0(73) & in_0(41) & in_0(9) & in_1(233) & in_1(201) & in_1(169) & in_1(137) & in_1(105);
mux_input_106 <= in_0(74) & in_0(42) & in_0(10) & in_1(234) & in_1(202) & in_1(170) & in_1(138) & in_1(106);
mux_input_107 <= in_0(75) & in_0(43) & in_0(11) & in_1(235) & in_1(203) & in_1(171) & in_1(139) & in_1(107);
mux_input_108 <= in_0(76) & in_0(44) & in_0(12) & in_1(236) & in_1(204) & in_1(172) & in_1(140) & in_1(108);
mux_input_109 <= in_0(77) & in_0(45) & in_0(13) & in_1(237) & in_1(205) & in_1(173) & in_1(141) & in_1(109);
mux_input_110 <= in_0(78) & in_0(46) & in_0(14) & in_1(238) & in_1(206) & in_1(174) & in_1(142) & in_1(110);
mux_input_111 <= in_0(79) & in_0(47) & in_0(15) & in_1(239) & in_1(207) & in_1(175) & in_1(143) & in_1(111);
mux_input_112 <= in_0(80) & in_0(48) & in_0(16) & in_1(240) & in_1(208) & in_1(176) & in_1(144) & in_1(112);
mux_input_113 <= in_0(81) & in_0(49) & in_0(17) & in_1(241) & in_1(209) & in_1(177) & in_1(145) & in_1(113);
mux_input_114 <= in_0(82) & in_0(50) & in_0(18) & in_1(242) & in_1(210) & in_1(178) & in_1(146) & in_1(114);
mux_input_115 <= in_0(83) & in_0(51) & in_0(19) & in_1(243) & in_1(211) & in_1(179) & in_1(147) & in_1(115);
mux_input_116 <= in_0(84) & in_0(52) & in_0(20) & in_1(244) & in_1(212) & in_1(180) & in_1(148) & in_1(116);
mux_input_117 <= in_0(85) & in_0(53) & in_0(21) & in_1(245) & in_1(213) & in_1(181) & in_1(149) & in_1(117);
mux_input_118 <= in_0(86) & in_0(54) & in_0(22) & in_1(246) & in_1(214) & in_1(182) & in_1(150) & in_1(118);
mux_input_119 <= in_0(87) & in_0(55) & in_0(23) & in_1(247) & in_1(215) & in_1(183) & in_1(151) & in_1(119);
mux_input_120 <= in_0(88) & in_0(56) & in_0(24) & in_1(248) & in_1(216) & in_1(184) & in_1(152) & in_1(120);
mux_input_121 <= in_0(89) & in_0(57) & in_0(25) & in_1(249) & in_1(217) & in_1(185) & in_1(153) & in_1(121);
mux_input_122 <= in_0(90) & in_0(58) & in_0(26) & in_1(250) & in_1(218) & in_1(186) & in_1(154) & in_1(122);
mux_input_123 <= in_0(91) & in_0(59) & in_0(27) & in_1(251) & in_1(219) & in_1(187) & in_1(155) & in_1(123);
mux_input_124 <= in_0(92) & in_0(60) & in_0(28) & in_1(252) & in_1(220) & in_1(188) & in_1(156) & in_1(124);
mux_input_125 <= in_0(93) & in_0(61) & in_0(29) & in_1(253) & in_1(221) & in_1(189) & in_1(157) & in_1(125);
mux_input_126 <= in_0(94) & in_0(62) & in_0(30) & in_1(254) & in_1(222) & in_1(190) & in_1(158) & in_1(126);
mux_input_127 <= in_0(95) & in_0(63) & in_0(31) & in_1(255) & in_1(223) & in_1(191) & in_1(159) & in_1(127);
-- Muxes from 128 to 159:
mux_input_128 <= in_0(128) & in_0(64) & in_0(32) & in_0(0) & in_1(224) & in_1(192) & in_1(160) & in_1(128);
mux_input_129 <= in_0(129) & in_0(65) & in_0(33) & in_0(1) & in_1(225) & in_1(193) & in_1(161) & in_1(129);
mux_input_130 <= in_0(130) & in_0(66) & in_0(34) & in_0(2) & in_1(226) & in_1(194) & in_1(162) & in_1(130);
mux_input_131 <= in_0(131) & in_0(67) & in_0(35) & in_0(3) & in_1(227) & in_1(195) & in_1(163) & in_1(131);
mux_input_132 <= in_0(132) & in_0(68) & in_0(36) & in_0(4) & in_1(228) & in_1(196) & in_1(164) & in_1(132);
mux_input_133 <= in_0(133) & in_0(69) & in_0(37) & in_0(5) & in_1(229) & in_1(197) & in_1(165) & in_1(133);
mux_input_134 <= in_0(134) & in_0(70) & in_0(38) & in_0(6) & in_1(230) & in_1(198) & in_1(166) & in_1(134);
mux_input_135 <= in_0(135) & in_0(71) & in_0(39) & in_0(7) & in_1(231) & in_1(199) & in_1(167) & in_1(135);
mux_input_136 <= in_0(136) & in_0(72) & in_0(40) & in_0(8) & in_1(232) & in_1(200) & in_1(168) & in_1(136);
mux_input_137 <= in_0(137) & in_0(73) & in_0(41) & in_0(9) & in_1(233) & in_1(201) & in_1(169) & in_1(137);
mux_input_138 <= in_0(138) & in_0(74) & in_0(42) & in_0(10) & in_1(234) & in_1(202) & in_1(170) & in_1(138);
mux_input_139 <= in_0(139) & in_0(75) & in_0(43) & in_0(11) & in_1(235) & in_1(203) & in_1(171) & in_1(139);
mux_input_140 <= in_0(140) & in_0(76) & in_0(44) & in_0(12) & in_1(236) & in_1(204) & in_1(172) & in_1(140);
mux_input_141 <= in_0(141) & in_0(77) & in_0(45) & in_0(13) & in_1(237) & in_1(205) & in_1(173) & in_1(141);
mux_input_142 <= in_0(142) & in_0(78) & in_0(46) & in_0(14) & in_1(238) & in_1(206) & in_1(174) & in_1(142);
mux_input_143 <= in_0(143) & in_0(79) & in_0(47) & in_0(15) & in_1(239) & in_1(207) & in_1(175) & in_1(143);
mux_input_144 <= in_0(144) & in_0(80) & in_0(48) & in_0(16) & in_1(240) & in_1(208) & in_1(176) & in_1(144);
mux_input_145 <= in_0(145) & in_0(81) & in_0(49) & in_0(17) & in_1(241) & in_1(209) & in_1(177) & in_1(145);
mux_input_146 <= in_0(146) & in_0(82) & in_0(50) & in_0(18) & in_1(242) & in_1(210) & in_1(178) & in_1(146);
mux_input_147 <= in_0(147) & in_0(83) & in_0(51) & in_0(19) & in_1(243) & in_1(211) & in_1(179) & in_1(147);
mux_input_148 <= in_0(148) & in_0(84) & in_0(52) & in_0(20) & in_1(244) & in_1(212) & in_1(180) & in_1(148);
mux_input_149 <= in_0(149) & in_0(85) & in_0(53) & in_0(21) & in_1(245) & in_1(213) & in_1(181) & in_1(149);
mux_input_150 <= in_0(150) & in_0(86) & in_0(54) & in_0(22) & in_1(246) & in_1(214) & in_1(182) & in_1(150);
mux_input_151 <= in_0(151) & in_0(87) & in_0(55) & in_0(23) & in_1(247) & in_1(215) & in_1(183) & in_1(151);
mux_input_152 <= in_0(152) & in_0(88) & in_0(56) & in_0(24) & in_1(248) & in_1(216) & in_1(184) & in_1(152);
mux_input_153 <= in_0(153) & in_0(89) & in_0(57) & in_0(25) & in_1(249) & in_1(217) & in_1(185) & in_1(153);
mux_input_154 <= in_0(154) & in_0(90) & in_0(58) & in_0(26) & in_1(250) & in_1(218) & in_1(186) & in_1(154);
mux_input_155 <= in_0(155) & in_0(91) & in_0(59) & in_0(27) & in_1(251) & in_1(219) & in_1(187) & in_1(155);
mux_input_156 <= in_0(156) & in_0(92) & in_0(60) & in_0(28) & in_1(252) & in_1(220) & in_1(188) & in_1(156);
mux_input_157 <= in_0(157) & in_0(93) & in_0(61) & in_0(29) & in_1(253) & in_1(221) & in_1(189) & in_1(157);
mux_input_158 <= in_0(158) & in_0(94) & in_0(62) & in_0(30) & in_1(254) & in_1(222) & in_1(190) & in_1(158);
mux_input_159 <= in_0(159) & in_0(95) & in_0(63) & in_0(31) & in_1(255) & in_1(223) & in_1(191) & in_1(159);
-- Muxes from 160 to 191:
mux_input_160 <= in_0(128) & in_0(96) & in_0(64) & in_0(32) & in_0(0) & in_1(224) & in_1(192) & in_1(160);
mux_input_161 <= in_0(129) & in_0(97) & in_0(65) & in_0(33) & in_0(1) & in_1(225) & in_1(193) & in_1(161);
mux_input_162 <= in_0(130) & in_0(98) & in_0(66) & in_0(34) & in_0(2) & in_1(226) & in_1(194) & in_1(162);
mux_input_163 <= in_0(131) & in_0(99) & in_0(67) & in_0(35) & in_0(3) & in_1(227) & in_1(195) & in_1(163);
mux_input_164 <= in_0(132) & in_0(100) & in_0(68) & in_0(36) & in_0(4) & in_1(228) & in_1(196) & in_1(164);
mux_input_165 <= in_0(133) & in_0(101) & in_0(69) & in_0(37) & in_0(5) & in_1(229) & in_1(197) & in_1(165);
mux_input_166 <= in_0(134) & in_0(102) & in_0(70) & in_0(38) & in_0(6) & in_1(230) & in_1(198) & in_1(166);
mux_input_167 <= in_0(135) & in_0(103) & in_0(71) & in_0(39) & in_0(7) & in_1(231) & in_1(199) & in_1(167);
mux_input_168 <= in_0(136) & in_0(104) & in_0(72) & in_0(40) & in_0(8) & in_1(232) & in_1(200) & in_1(168);
mux_input_169 <= in_0(137) & in_0(105) & in_0(73) & in_0(41) & in_0(9) & in_1(233) & in_1(201) & in_1(169);
mux_input_170 <= in_0(138) & in_0(106) & in_0(74) & in_0(42) & in_0(10) & in_1(234) & in_1(202) & in_1(170);
mux_input_171 <= in_0(139) & in_0(107) & in_0(75) & in_0(43) & in_0(11) & in_1(235) & in_1(203) & in_1(171);
mux_input_172 <= in_0(140) & in_0(108) & in_0(76) & in_0(44) & in_0(12) & in_1(236) & in_1(204) & in_1(172);
mux_input_173 <= in_0(141) & in_0(109) & in_0(77) & in_0(45) & in_0(13) & in_1(237) & in_1(205) & in_1(173);
mux_input_174 <= in_0(142) & in_0(110) & in_0(78) & in_0(46) & in_0(14) & in_1(238) & in_1(206) & in_1(174);
mux_input_175 <= in_0(143) & in_0(111) & in_0(79) & in_0(47) & in_0(15) & in_1(239) & in_1(207) & in_1(175);
mux_input_176 <= in_0(144) & in_0(112) & in_0(80) & in_0(48) & in_0(16) & in_1(240) & in_1(208) & in_1(176);
mux_input_177 <= in_0(145) & in_0(113) & in_0(81) & in_0(49) & in_0(17) & in_1(241) & in_1(209) & in_1(177);
mux_input_178 <= in_0(146) & in_0(114) & in_0(82) & in_0(50) & in_0(18) & in_1(242) & in_1(210) & in_1(178);
mux_input_179 <= in_0(147) & in_0(115) & in_0(83) & in_0(51) & in_0(19) & in_1(243) & in_1(211) & in_1(179);
mux_input_180 <= in_0(148) & in_0(116) & in_0(84) & in_0(52) & in_0(20) & in_1(244) & in_1(212) & in_1(180);
mux_input_181 <= in_0(149) & in_0(117) & in_0(85) & in_0(53) & in_0(21) & in_1(245) & in_1(213) & in_1(181);
mux_input_182 <= in_0(150) & in_0(118) & in_0(86) & in_0(54) & in_0(22) & in_1(246) & in_1(214) & in_1(182);
mux_input_183 <= in_0(151) & in_0(119) & in_0(87) & in_0(55) & in_0(23) & in_1(247) & in_1(215) & in_1(183);
mux_input_184 <= in_0(152) & in_0(120) & in_0(88) & in_0(56) & in_0(24) & in_1(248) & in_1(216) & in_1(184);
mux_input_185 <= in_0(153) & in_0(121) & in_0(89) & in_0(57) & in_0(25) & in_1(249) & in_1(217) & in_1(185);
mux_input_186 <= in_0(154) & in_0(122) & in_0(90) & in_0(58) & in_0(26) & in_1(250) & in_1(218) & in_1(186);
mux_input_187 <= in_0(155) & in_0(123) & in_0(91) & in_0(59) & in_0(27) & in_1(251) & in_1(219) & in_1(187);
mux_input_188 <= in_0(156) & in_0(124) & in_0(92) & in_0(60) & in_0(28) & in_1(252) & in_1(220) & in_1(188);
mux_input_189 <= in_0(157) & in_0(125) & in_0(93) & in_0(61) & in_0(29) & in_1(253) & in_1(221) & in_1(189);
mux_input_190 <= in_0(158) & in_0(126) & in_0(94) & in_0(62) & in_0(30) & in_1(254) & in_1(222) & in_1(190);
mux_input_191 <= in_0(159) & in_0(127) & in_0(95) & in_0(63) & in_0(31) & in_1(255) & in_1(223) & in_1(191);
-- Muxes from 192 to 223:
mux_input_192 <= in_0(160) & in_0(128) & in_0(96) & in_0(64) & in_0(32) & in_0(0) & in_1(224) & in_1(192);
mux_input_193 <= in_0(161) & in_0(129) & in_0(97) & in_0(65) & in_0(33) & in_0(1) & in_1(225) & in_1(193);
mux_input_194 <= in_0(162) & in_0(130) & in_0(98) & in_0(66) & in_0(34) & in_0(2) & in_1(226) & in_1(194);
mux_input_195 <= in_0(163) & in_0(131) & in_0(99) & in_0(67) & in_0(35) & in_0(3) & in_1(227) & in_1(195);
mux_input_196 <= in_0(164) & in_0(132) & in_0(100) & in_0(68) & in_0(36) & in_0(4) & in_1(228) & in_1(196);
mux_input_197 <= in_0(165) & in_0(133) & in_0(101) & in_0(69) & in_0(37) & in_0(5) & in_1(229) & in_1(197);
mux_input_198 <= in_0(166) & in_0(134) & in_0(102) & in_0(70) & in_0(38) & in_0(6) & in_1(230) & in_1(198);
mux_input_199 <= in_0(167) & in_0(135) & in_0(103) & in_0(71) & in_0(39) & in_0(7) & in_1(231) & in_1(199);
mux_input_200 <= in_0(168) & in_0(136) & in_0(104) & in_0(72) & in_0(40) & in_0(8) & in_1(232) & in_1(200);
mux_input_201 <= in_0(169) & in_0(137) & in_0(105) & in_0(73) & in_0(41) & in_0(9) & in_1(233) & in_1(201);
mux_input_202 <= in_0(170) & in_0(138) & in_0(106) & in_0(74) & in_0(42) & in_0(10) & in_1(234) & in_1(202);
mux_input_203 <= in_0(171) & in_0(139) & in_0(107) & in_0(75) & in_0(43) & in_0(11) & in_1(235) & in_1(203);
mux_input_204 <= in_0(172) & in_0(140) & in_0(108) & in_0(76) & in_0(44) & in_0(12) & in_1(236) & in_1(204);
mux_input_205 <= in_0(173) & in_0(141) & in_0(109) & in_0(77) & in_0(45) & in_0(13) & in_1(237) & in_1(205);
mux_input_206 <= in_0(174) & in_0(142) & in_0(110) & in_0(78) & in_0(46) & in_0(14) & in_1(238) & in_1(206);
mux_input_207 <= in_0(175) & in_0(143) & in_0(111) & in_0(79) & in_0(47) & in_0(15) & in_1(239) & in_1(207);
mux_input_208 <= in_0(176) & in_0(144) & in_0(112) & in_0(80) & in_0(48) & in_0(16) & in_1(240) & in_1(208);
mux_input_209 <= in_0(177) & in_0(145) & in_0(113) & in_0(81) & in_0(49) & in_0(17) & in_1(241) & in_1(209);
mux_input_210 <= in_0(178) & in_0(146) & in_0(114) & in_0(82) & in_0(50) & in_0(18) & in_1(242) & in_1(210);
mux_input_211 <= in_0(179) & in_0(147) & in_0(115) & in_0(83) & in_0(51) & in_0(19) & in_1(243) & in_1(211);
mux_input_212 <= in_0(180) & in_0(148) & in_0(116) & in_0(84) & in_0(52) & in_0(20) & in_1(244) & in_1(212);
mux_input_213 <= in_0(181) & in_0(149) & in_0(117) & in_0(85) & in_0(53) & in_0(21) & in_1(245) & in_1(213);
mux_input_214 <= in_0(182) & in_0(150) & in_0(118) & in_0(86) & in_0(54) & in_0(22) & in_1(246) & in_1(214);
mux_input_215 <= in_0(183) & in_0(151) & in_0(119) & in_0(87) & in_0(55) & in_0(23) & in_1(247) & in_1(215);
mux_input_216 <= in_0(184) & in_0(152) & in_0(120) & in_0(88) & in_0(56) & in_0(24) & in_1(248) & in_1(216);
mux_input_217 <= in_0(185) & in_0(153) & in_0(121) & in_0(89) & in_0(57) & in_0(25) & in_1(249) & in_1(217);
mux_input_218 <= in_0(186) & in_0(154) & in_0(122) & in_0(90) & in_0(58) & in_0(26) & in_1(250) & in_1(218);
mux_input_219 <= in_0(187) & in_0(155) & in_0(123) & in_0(91) & in_0(59) & in_0(27) & in_1(251) & in_1(219);
mux_input_220 <= in_0(188) & in_0(156) & in_0(124) & in_0(92) & in_0(60) & in_0(28) & in_1(252) & in_1(220);
mux_input_221 <= in_0(189) & in_0(157) & in_0(125) & in_0(93) & in_0(61) & in_0(29) & in_1(253) & in_1(221);
mux_input_222 <= in_0(190) & in_0(158) & in_0(126) & in_0(94) & in_0(62) & in_0(30) & in_1(254) & in_1(222);
mux_input_223 <= in_0(191) & in_0(159) & in_0(127) & in_0(95) & in_0(63) & in_0(31) & in_1(255) & in_1(223);
-- Muxes from 224 to 255:
mux_input_224 <= in_0(192) & in_0(160) & in_0(128) & in_0(96) & in_0(64) & in_0(32) & in_0(0) & in_1(224);
mux_input_225 <= in_0(193) & in_0(161) & in_0(129) & in_0(97) & in_0(65) & in_0(33) & in_0(1) & in_1(225);
mux_input_226 <= in_0(194) & in_0(162) & in_0(130) & in_0(98) & in_0(66) & in_0(34) & in_0(2) & in_1(226);
mux_input_227 <= in_0(195) & in_0(163) & in_0(131) & in_0(99) & in_0(67) & in_0(35) & in_0(3) & in_1(227);
mux_input_228 <= in_0(196) & in_0(164) & in_0(132) & in_0(100) & in_0(68) & in_0(36) & in_0(4) & in_1(228);
mux_input_229 <= in_0(197) & in_0(165) & in_0(133) & in_0(101) & in_0(69) & in_0(37) & in_0(5) & in_1(229);
mux_input_230 <= in_0(198) & in_0(166) & in_0(134) & in_0(102) & in_0(70) & in_0(38) & in_0(6) & in_1(230);
mux_input_231 <= in_0(199) & in_0(167) & in_0(135) & in_0(103) & in_0(71) & in_0(39) & in_0(7) & in_1(231);
mux_input_232 <= in_0(200) & in_0(168) & in_0(136) & in_0(104) & in_0(72) & in_0(40) & in_0(8) & in_1(232);
mux_input_233 <= in_0(201) & in_0(169) & in_0(137) & in_0(105) & in_0(73) & in_0(41) & in_0(9) & in_1(233);
mux_input_234 <= in_0(202) & in_0(170) & in_0(138) & in_0(106) & in_0(74) & in_0(42) & in_0(10) & in_1(234);
mux_input_235 <= in_0(203) & in_0(171) & in_0(139) & in_0(107) & in_0(75) & in_0(43) & in_0(11) & in_1(235);
mux_input_236 <= in_0(204) & in_0(172) & in_0(140) & in_0(108) & in_0(76) & in_0(44) & in_0(12) & in_1(236);
mux_input_237 <= in_0(205) & in_0(173) & in_0(141) & in_0(109) & in_0(77) & in_0(45) & in_0(13) & in_1(237);
mux_input_238 <= in_0(206) & in_0(174) & in_0(142) & in_0(110) & in_0(78) & in_0(46) & in_0(14) & in_1(238);
mux_input_239 <= in_0(207) & in_0(175) & in_0(143) & in_0(111) & in_0(79) & in_0(47) & in_0(15) & in_1(239);
mux_input_240 <= in_0(208) & in_0(176) & in_0(144) & in_0(112) & in_0(80) & in_0(48) & in_0(16) & in_1(240);
mux_input_241 <= in_0(209) & in_0(177) & in_0(145) & in_0(113) & in_0(81) & in_0(49) & in_0(17) & in_1(241);
mux_input_242 <= in_0(210) & in_0(178) & in_0(146) & in_0(114) & in_0(82) & in_0(50) & in_0(18) & in_1(242);
mux_input_243 <= in_0(211) & in_0(179) & in_0(147) & in_0(115) & in_0(83) & in_0(51) & in_0(19) & in_1(243);
mux_input_244 <= in_0(212) & in_0(180) & in_0(148) & in_0(116) & in_0(84) & in_0(52) & in_0(20) & in_1(244);
mux_input_245 <= in_0(213) & in_0(181) & in_0(149) & in_0(117) & in_0(85) & in_0(53) & in_0(21) & in_1(245);
mux_input_246 <= in_0(214) & in_0(182) & in_0(150) & in_0(118) & in_0(86) & in_0(54) & in_0(22) & in_1(246);
mux_input_247 <= in_0(215) & in_0(183) & in_0(151) & in_0(119) & in_0(87) & in_0(55) & in_0(23) & in_1(247);
mux_input_248 <= in_0(216) & in_0(184) & in_0(152) & in_0(120) & in_0(88) & in_0(56) & in_0(24) & in_1(248);
mux_input_249 <= in_0(217) & in_0(185) & in_0(153) & in_0(121) & in_0(89) & in_0(57) & in_0(25) & in_1(249);
mux_input_250 <= in_0(218) & in_0(186) & in_0(154) & in_0(122) & in_0(90) & in_0(58) & in_0(26) & in_1(250);
mux_input_251 <= in_0(219) & in_0(187) & in_0(155) & in_0(123) & in_0(91) & in_0(59) & in_0(27) & in_1(251);
mux_input_252 <= in_0(220) & in_0(188) & in_0(156) & in_0(124) & in_0(92) & in_0(60) & in_0(28) & in_1(252);
mux_input_253 <= in_0(221) & in_0(189) & in_0(157) & in_0(125) & in_0(93) & in_0(61) & in_0(29) & in_1(253);
mux_input_254 <= in_0(222) & in_0(190) & in_0(158) & in_0(126) & in_0(94) & in_0(62) & in_0(30) & in_1(254);
mux_input_255 <= in_0(223) & in_0(191) & in_0(159) & in_0(127) & in_0(95) & in_0(63) & in_0(31) & in_1(255);
-- Port maps:
inst_mux_0: entity work.mux8 port map(mux_input_0, sel_mux, data_out(0));
inst_mux_1: entity work.mux8 port map(mux_input_1, sel_mux, data_out(1));
inst_mux_2: entity work.mux8 port map(mux_input_2, sel_mux, data_out(2));
inst_mux_3: entity work.mux8 port map(mux_input_3, sel_mux, data_out(3));
inst_mux_4: entity work.mux8 port map(mux_input_4, sel_mux, data_out(4));
inst_mux_5: entity work.mux8 port map(mux_input_5, sel_mux, data_out(5));
inst_mux_6: entity work.mux8 port map(mux_input_6, sel_mux, data_out(6));
inst_mux_7: entity work.mux8 port map(mux_input_7, sel_mux, data_out(7));
inst_mux_8: entity work.mux8 port map(mux_input_8, sel_mux, data_out(8));
inst_mux_9: entity work.mux8 port map(mux_input_9, sel_mux, data_out(9));
inst_mux_10: entity work.mux8 port map(mux_input_10, sel_mux, data_out(10));
inst_mux_11: entity work.mux8 port map(mux_input_11, sel_mux, data_out(11));
inst_mux_12: entity work.mux8 port map(mux_input_12, sel_mux, data_out(12));
inst_mux_13: entity work.mux8 port map(mux_input_13, sel_mux, data_out(13));
inst_mux_14: entity work.mux8 port map(mux_input_14, sel_mux, data_out(14));
inst_mux_15: entity work.mux8 port map(mux_input_15, sel_mux, data_out(15));
inst_mux_16: entity work.mux8 port map(mux_input_16, sel_mux, data_out(16));
inst_mux_17: entity work.mux8 port map(mux_input_17, sel_mux, data_out(17));
inst_mux_18: entity work.mux8 port map(mux_input_18, sel_mux, data_out(18));
inst_mux_19: entity work.mux8 port map(mux_input_19, sel_mux, data_out(19));
inst_mux_20: entity work.mux8 port map(mux_input_20, sel_mux, data_out(20));
inst_mux_21: entity work.mux8 port map(mux_input_21, sel_mux, data_out(21));
inst_mux_22: entity work.mux8 port map(mux_input_22, sel_mux, data_out(22));
inst_mux_23: entity work.mux8 port map(mux_input_23, sel_mux, data_out(23));
inst_mux_24: entity work.mux8 port map(mux_input_24, sel_mux, data_out(24));
inst_mux_25: entity work.mux8 port map(mux_input_25, sel_mux, data_out(25));
inst_mux_26: entity work.mux8 port map(mux_input_26, sel_mux, data_out(26));
inst_mux_27: entity work.mux8 port map(mux_input_27, sel_mux, data_out(27));
inst_mux_28: entity work.mux8 port map(mux_input_28, sel_mux, data_out(28));
inst_mux_29: entity work.mux8 port map(mux_input_29, sel_mux, data_out(29));
inst_mux_30: entity work.mux8 port map(mux_input_30, sel_mux, data_out(30));
inst_mux_31: entity work.mux8 port map(mux_input_31, sel_mux, data_out(31));
inst_mux_32: entity work.mux8 port map(mux_input_32, sel_mux, data_out(32));
inst_mux_33: entity work.mux8 port map(mux_input_33, sel_mux, data_out(33));
inst_mux_34: entity work.mux8 port map(mux_input_34, sel_mux, data_out(34));
inst_mux_35: entity work.mux8 port map(mux_input_35, sel_mux, data_out(35));
inst_mux_36: entity work.mux8 port map(mux_input_36, sel_mux, data_out(36));
inst_mux_37: entity work.mux8 port map(mux_input_37, sel_mux, data_out(37));
inst_mux_38: entity work.mux8 port map(mux_input_38, sel_mux, data_out(38));
inst_mux_39: entity work.mux8 port map(mux_input_39, sel_mux, data_out(39));
inst_mux_40: entity work.mux8 port map(mux_input_40, sel_mux, data_out(40));
inst_mux_41: entity work.mux8 port map(mux_input_41, sel_mux, data_out(41));
inst_mux_42: entity work.mux8 port map(mux_input_42, sel_mux, data_out(42));
inst_mux_43: entity work.mux8 port map(mux_input_43, sel_mux, data_out(43));
inst_mux_44: entity work.mux8 port map(mux_input_44, sel_mux, data_out(44));
inst_mux_45: entity work.mux8 port map(mux_input_45, sel_mux, data_out(45));
inst_mux_46: entity work.mux8 port map(mux_input_46, sel_mux, data_out(46));
inst_mux_47: entity work.mux8 port map(mux_input_47, sel_mux, data_out(47));
inst_mux_48: entity work.mux8 port map(mux_input_48, sel_mux, data_out(48));
inst_mux_49: entity work.mux8 port map(mux_input_49, sel_mux, data_out(49));
inst_mux_50: entity work.mux8 port map(mux_input_50, sel_mux, data_out(50));
inst_mux_51: entity work.mux8 port map(mux_input_51, sel_mux, data_out(51));
inst_mux_52: entity work.mux8 port map(mux_input_52, sel_mux, data_out(52));
inst_mux_53: entity work.mux8 port map(mux_input_53, sel_mux, data_out(53));
inst_mux_54: entity work.mux8 port map(mux_input_54, sel_mux, data_out(54));
inst_mux_55: entity work.mux8 port map(mux_input_55, sel_mux, data_out(55));
inst_mux_56: entity work.mux8 port map(mux_input_56, sel_mux, data_out(56));
inst_mux_57: entity work.mux8 port map(mux_input_57, sel_mux, data_out(57));
inst_mux_58: entity work.mux8 port map(mux_input_58, sel_mux, data_out(58));
inst_mux_59: entity work.mux8 port map(mux_input_59, sel_mux, data_out(59));
inst_mux_60: entity work.mux8 port map(mux_input_60, sel_mux, data_out(60));
inst_mux_61: entity work.mux8 port map(mux_input_61, sel_mux, data_out(61));
inst_mux_62: entity work.mux8 port map(mux_input_62, sel_mux, data_out(62));
inst_mux_63: entity work.mux8 port map(mux_input_63, sel_mux, data_out(63));
inst_mux_64: entity work.mux8 port map(mux_input_64, sel_mux, data_out(64));
inst_mux_65: entity work.mux8 port map(mux_input_65, sel_mux, data_out(65));
inst_mux_66: entity work.mux8 port map(mux_input_66, sel_mux, data_out(66));
inst_mux_67: entity work.mux8 port map(mux_input_67, sel_mux, data_out(67));
inst_mux_68: entity work.mux8 port map(mux_input_68, sel_mux, data_out(68));
inst_mux_69: entity work.mux8 port map(mux_input_69, sel_mux, data_out(69));
inst_mux_70: entity work.mux8 port map(mux_input_70, sel_mux, data_out(70));
inst_mux_71: entity work.mux8 port map(mux_input_71, sel_mux, data_out(71));
inst_mux_72: entity work.mux8 port map(mux_input_72, sel_mux, data_out(72));
inst_mux_73: entity work.mux8 port map(mux_input_73, sel_mux, data_out(73));
inst_mux_74: entity work.mux8 port map(mux_input_74, sel_mux, data_out(74));
inst_mux_75: entity work.mux8 port map(mux_input_75, sel_mux, data_out(75));
inst_mux_76: entity work.mux8 port map(mux_input_76, sel_mux, data_out(76));
inst_mux_77: entity work.mux8 port map(mux_input_77, sel_mux, data_out(77));
inst_mux_78: entity work.mux8 port map(mux_input_78, sel_mux, data_out(78));
inst_mux_79: entity work.mux8 port map(mux_input_79, sel_mux, data_out(79));
inst_mux_80: entity work.mux8 port map(mux_input_80, sel_mux, data_out(80));
inst_mux_81: entity work.mux8 port map(mux_input_81, sel_mux, data_out(81));
inst_mux_82: entity work.mux8 port map(mux_input_82, sel_mux, data_out(82));
inst_mux_83: entity work.mux8 port map(mux_input_83, sel_mux, data_out(83));
inst_mux_84: entity work.mux8 port map(mux_input_84, sel_mux, data_out(84));
inst_mux_85: entity work.mux8 port map(mux_input_85, sel_mux, data_out(85));
inst_mux_86: entity work.mux8 port map(mux_input_86, sel_mux, data_out(86));
inst_mux_87: entity work.mux8 port map(mux_input_87, sel_mux, data_out(87));
inst_mux_88: entity work.mux8 port map(mux_input_88, sel_mux, data_out(88));
inst_mux_89: entity work.mux8 port map(mux_input_89, sel_mux, data_out(89));
inst_mux_90: entity work.mux8 port map(mux_input_90, sel_mux, data_out(90));
inst_mux_91: entity work.mux8 port map(mux_input_91, sel_mux, data_out(91));
inst_mux_92: entity work.mux8 port map(mux_input_92, sel_mux, data_out(92));
inst_mux_93: entity work.mux8 port map(mux_input_93, sel_mux, data_out(93));
inst_mux_94: entity work.mux8 port map(mux_input_94, sel_mux, data_out(94));
inst_mux_95: entity work.mux8 port map(mux_input_95, sel_mux, data_out(95));
inst_mux_96: entity work.mux8 port map(mux_input_96, sel_mux, data_out(96));
inst_mux_97: entity work.mux8 port map(mux_input_97, sel_mux, data_out(97));
inst_mux_98: entity work.mux8 port map(mux_input_98, sel_mux, data_out(98));
inst_mux_99: entity work.mux8 port map(mux_input_99, sel_mux, data_out(99));
inst_mux_100: entity work.mux8 port map(mux_input_100, sel_mux, data_out(100));
inst_mux_101: entity work.mux8 port map(mux_input_101, sel_mux, data_out(101));
inst_mux_102: entity work.mux8 port map(mux_input_102, sel_mux, data_out(102));
inst_mux_103: entity work.mux8 port map(mux_input_103, sel_mux, data_out(103));
inst_mux_104: entity work.mux8 port map(mux_input_104, sel_mux, data_out(104));
inst_mux_105: entity work.mux8 port map(mux_input_105, sel_mux, data_out(105));
inst_mux_106: entity work.mux8 port map(mux_input_106, sel_mux, data_out(106));
inst_mux_107: entity work.mux8 port map(mux_input_107, sel_mux, data_out(107));
inst_mux_108: entity work.mux8 port map(mux_input_108, sel_mux, data_out(108));
inst_mux_109: entity work.mux8 port map(mux_input_109, sel_mux, data_out(109));
inst_mux_110: entity work.mux8 port map(mux_input_110, sel_mux, data_out(110));
inst_mux_111: entity work.mux8 port map(mux_input_111, sel_mux, data_out(111));
inst_mux_112: entity work.mux8 port map(mux_input_112, sel_mux, data_out(112));
inst_mux_113: entity work.mux8 port map(mux_input_113, sel_mux, data_out(113));
inst_mux_114: entity work.mux8 port map(mux_input_114, sel_mux, data_out(114));
inst_mux_115: entity work.mux8 port map(mux_input_115, sel_mux, data_out(115));
inst_mux_116: entity work.mux8 port map(mux_input_116, sel_mux, data_out(116));
inst_mux_117: entity work.mux8 port map(mux_input_117, sel_mux, data_out(117));
inst_mux_118: entity work.mux8 port map(mux_input_118, sel_mux, data_out(118));
inst_mux_119: entity work.mux8 port map(mux_input_119, sel_mux, data_out(119));
inst_mux_120: entity work.mux8 port map(mux_input_120, sel_mux, data_out(120));
inst_mux_121: entity work.mux8 port map(mux_input_121, sel_mux, data_out(121));
inst_mux_122: entity work.mux8 port map(mux_input_122, sel_mux, data_out(122));
inst_mux_123: entity work.mux8 port map(mux_input_123, sel_mux, data_out(123));
inst_mux_124: entity work.mux8 port map(mux_input_124, sel_mux, data_out(124));
inst_mux_125: entity work.mux8 port map(mux_input_125, sel_mux, data_out(125));
inst_mux_126: entity work.mux8 port map(mux_input_126, sel_mux, data_out(126));
inst_mux_127: entity work.mux8 port map(mux_input_127, sel_mux, data_out(127));
inst_mux_128: entity work.mux8 port map(mux_input_128, sel_mux, data_out(128));
inst_mux_129: entity work.mux8 port map(mux_input_129, sel_mux, data_out(129));
inst_mux_130: entity work.mux8 port map(mux_input_130, sel_mux, data_out(130));
inst_mux_131: entity work.mux8 port map(mux_input_131, sel_mux, data_out(131));
inst_mux_132: entity work.mux8 port map(mux_input_132, sel_mux, data_out(132));
inst_mux_133: entity work.mux8 port map(mux_input_133, sel_mux, data_out(133));
inst_mux_134: entity work.mux8 port map(mux_input_134, sel_mux, data_out(134));
inst_mux_135: entity work.mux8 port map(mux_input_135, sel_mux, data_out(135));
inst_mux_136: entity work.mux8 port map(mux_input_136, sel_mux, data_out(136));
inst_mux_137: entity work.mux8 port map(mux_input_137, sel_mux, data_out(137));
inst_mux_138: entity work.mux8 port map(mux_input_138, sel_mux, data_out(138));
inst_mux_139: entity work.mux8 port map(mux_input_139, sel_mux, data_out(139));
inst_mux_140: entity work.mux8 port map(mux_input_140, sel_mux, data_out(140));
inst_mux_141: entity work.mux8 port map(mux_input_141, sel_mux, data_out(141));
inst_mux_142: entity work.mux8 port map(mux_input_142, sel_mux, data_out(142));
inst_mux_143: entity work.mux8 port map(mux_input_143, sel_mux, data_out(143));
inst_mux_144: entity work.mux8 port map(mux_input_144, sel_mux, data_out(144));
inst_mux_145: entity work.mux8 port map(mux_input_145, sel_mux, data_out(145));
inst_mux_146: entity work.mux8 port map(mux_input_146, sel_mux, data_out(146));
inst_mux_147: entity work.mux8 port map(mux_input_147, sel_mux, data_out(147));
inst_mux_148: entity work.mux8 port map(mux_input_148, sel_mux, data_out(148));
inst_mux_149: entity work.mux8 port map(mux_input_149, sel_mux, data_out(149));
inst_mux_150: entity work.mux8 port map(mux_input_150, sel_mux, data_out(150));
inst_mux_151: entity work.mux8 port map(mux_input_151, sel_mux, data_out(151));
inst_mux_152: entity work.mux8 port map(mux_input_152, sel_mux, data_out(152));
inst_mux_153: entity work.mux8 port map(mux_input_153, sel_mux, data_out(153));
inst_mux_154: entity work.mux8 port map(mux_input_154, sel_mux, data_out(154));
inst_mux_155: entity work.mux8 port map(mux_input_155, sel_mux, data_out(155));
inst_mux_156: entity work.mux8 port map(mux_input_156, sel_mux, data_out(156));
inst_mux_157: entity work.mux8 port map(mux_input_157, sel_mux, data_out(157));
inst_mux_158: entity work.mux8 port map(mux_input_158, sel_mux, data_out(158));
inst_mux_159: entity work.mux8 port map(mux_input_159, sel_mux, data_out(159));
inst_mux_160: entity work.mux8 port map(mux_input_160, sel_mux, data_out(160));
inst_mux_161: entity work.mux8 port map(mux_input_161, sel_mux, data_out(161));
inst_mux_162: entity work.mux8 port map(mux_input_162, sel_mux, data_out(162));
inst_mux_163: entity work.mux8 port map(mux_input_163, sel_mux, data_out(163));
inst_mux_164: entity work.mux8 port map(mux_input_164, sel_mux, data_out(164));
inst_mux_165: entity work.mux8 port map(mux_input_165, sel_mux, data_out(165));
inst_mux_166: entity work.mux8 port map(mux_input_166, sel_mux, data_out(166));
inst_mux_167: entity work.mux8 port map(mux_input_167, sel_mux, data_out(167));
inst_mux_168: entity work.mux8 port map(mux_input_168, sel_mux, data_out(168));
inst_mux_169: entity work.mux8 port map(mux_input_169, sel_mux, data_out(169));
inst_mux_170: entity work.mux8 port map(mux_input_170, sel_mux, data_out(170));
inst_mux_171: entity work.mux8 port map(mux_input_171, sel_mux, data_out(171));
inst_mux_172: entity work.mux8 port map(mux_input_172, sel_mux, data_out(172));
inst_mux_173: entity work.mux8 port map(mux_input_173, sel_mux, data_out(173));
inst_mux_174: entity work.mux8 port map(mux_input_174, sel_mux, data_out(174));
inst_mux_175: entity work.mux8 port map(mux_input_175, sel_mux, data_out(175));
inst_mux_176: entity work.mux8 port map(mux_input_176, sel_mux, data_out(176));
inst_mux_177: entity work.mux8 port map(mux_input_177, sel_mux, data_out(177));
inst_mux_178: entity work.mux8 port map(mux_input_178, sel_mux, data_out(178));
inst_mux_179: entity work.mux8 port map(mux_input_179, sel_mux, data_out(179));
inst_mux_180: entity work.mux8 port map(mux_input_180, sel_mux, data_out(180));
inst_mux_181: entity work.mux8 port map(mux_input_181, sel_mux, data_out(181));
inst_mux_182: entity work.mux8 port map(mux_input_182, sel_mux, data_out(182));
inst_mux_183: entity work.mux8 port map(mux_input_183, sel_mux, data_out(183));
inst_mux_184: entity work.mux8 port map(mux_input_184, sel_mux, data_out(184));
inst_mux_185: entity work.mux8 port map(mux_input_185, sel_mux, data_out(185));
inst_mux_186: entity work.mux8 port map(mux_input_186, sel_mux, data_out(186));
inst_mux_187: entity work.mux8 port map(mux_input_187, sel_mux, data_out(187));
inst_mux_188: entity work.mux8 port map(mux_input_188, sel_mux, data_out(188));
inst_mux_189: entity work.mux8 port map(mux_input_189, sel_mux, data_out(189));
inst_mux_190: entity work.mux8 port map(mux_input_190, sel_mux, data_out(190));
inst_mux_191: entity work.mux8 port map(mux_input_191, sel_mux, data_out(191));
inst_mux_192: entity work.mux8 port map(mux_input_192, sel_mux, data_out(192));
inst_mux_193: entity work.mux8 port map(mux_input_193, sel_mux, data_out(193));
inst_mux_194: entity work.mux8 port map(mux_input_194, sel_mux, data_out(194));
inst_mux_195: entity work.mux8 port map(mux_input_195, sel_mux, data_out(195));
inst_mux_196: entity work.mux8 port map(mux_input_196, sel_mux, data_out(196));
inst_mux_197: entity work.mux8 port map(mux_input_197, sel_mux, data_out(197));
inst_mux_198: entity work.mux8 port map(mux_input_198, sel_mux, data_out(198));
inst_mux_199: entity work.mux8 port map(mux_input_199, sel_mux, data_out(199));
inst_mux_200: entity work.mux8 port map(mux_input_200, sel_mux, data_out(200));
inst_mux_201: entity work.mux8 port map(mux_input_201, sel_mux, data_out(201));
inst_mux_202: entity work.mux8 port map(mux_input_202, sel_mux, data_out(202));
inst_mux_203: entity work.mux8 port map(mux_input_203, sel_mux, data_out(203));
inst_mux_204: entity work.mux8 port map(mux_input_204, sel_mux, data_out(204));
inst_mux_205: entity work.mux8 port map(mux_input_205, sel_mux, data_out(205));
inst_mux_206: entity work.mux8 port map(mux_input_206, sel_mux, data_out(206));
inst_mux_207: entity work.mux8 port map(mux_input_207, sel_mux, data_out(207));
inst_mux_208: entity work.mux8 port map(mux_input_208, sel_mux, data_out(208));
inst_mux_209: entity work.mux8 port map(mux_input_209, sel_mux, data_out(209));
inst_mux_210: entity work.mux8 port map(mux_input_210, sel_mux, data_out(210));
inst_mux_211: entity work.mux8 port map(mux_input_211, sel_mux, data_out(211));
inst_mux_212: entity work.mux8 port map(mux_input_212, sel_mux, data_out(212));
inst_mux_213: entity work.mux8 port map(mux_input_213, sel_mux, data_out(213));
inst_mux_214: entity work.mux8 port map(mux_input_214, sel_mux, data_out(214));
inst_mux_215: entity work.mux8 port map(mux_input_215, sel_mux, data_out(215));
inst_mux_216: entity work.mux8 port map(mux_input_216, sel_mux, data_out(216));
inst_mux_217: entity work.mux8 port map(mux_input_217, sel_mux, data_out(217));
inst_mux_218: entity work.mux8 port map(mux_input_218, sel_mux, data_out(218));
inst_mux_219: entity work.mux8 port map(mux_input_219, sel_mux, data_out(219));
inst_mux_220: entity work.mux8 port map(mux_input_220, sel_mux, data_out(220));
inst_mux_221: entity work.mux8 port map(mux_input_221, sel_mux, data_out(221));
inst_mux_222: entity work.mux8 port map(mux_input_222, sel_mux, data_out(222));
inst_mux_223: entity work.mux8 port map(mux_input_223, sel_mux, data_out(223));
inst_mux_224: entity work.mux8 port map(mux_input_224, sel_mux, data_out(224));
inst_mux_225: entity work.mux8 port map(mux_input_225, sel_mux, data_out(225));
inst_mux_226: entity work.mux8 port map(mux_input_226, sel_mux, data_out(226));
inst_mux_227: entity work.mux8 port map(mux_input_227, sel_mux, data_out(227));
inst_mux_228: entity work.mux8 port map(mux_input_228, sel_mux, data_out(228));
inst_mux_229: entity work.mux8 port map(mux_input_229, sel_mux, data_out(229));
inst_mux_230: entity work.mux8 port map(mux_input_230, sel_mux, data_out(230));
inst_mux_231: entity work.mux8 port map(mux_input_231, sel_mux, data_out(231));
inst_mux_232: entity work.mux8 port map(mux_input_232, sel_mux, data_out(232));
inst_mux_233: entity work.mux8 port map(mux_input_233, sel_mux, data_out(233));
inst_mux_234: entity work.mux8 port map(mux_input_234, sel_mux, data_out(234));
inst_mux_235: entity work.mux8 port map(mux_input_235, sel_mux, data_out(235));
inst_mux_236: entity work.mux8 port map(mux_input_236, sel_mux, data_out(236));
inst_mux_237: entity work.mux8 port map(mux_input_237, sel_mux, data_out(237));
inst_mux_238: entity work.mux8 port map(mux_input_238, sel_mux, data_out(238));
inst_mux_239: entity work.mux8 port map(mux_input_239, sel_mux, data_out(239));
inst_mux_240: entity work.mux8 port map(mux_input_240, sel_mux, data_out(240));
inst_mux_241: entity work.mux8 port map(mux_input_241, sel_mux, data_out(241));
inst_mux_242: entity work.mux8 port map(mux_input_242, sel_mux, data_out(242));
inst_mux_243: entity work.mux8 port map(mux_input_243, sel_mux, data_out(243));
inst_mux_244: entity work.mux8 port map(mux_input_244, sel_mux, data_out(244));
inst_mux_245: entity work.mux8 port map(mux_input_245, sel_mux, data_out(245));
inst_mux_246: entity work.mux8 port map(mux_input_246, sel_mux, data_out(246));
inst_mux_247: entity work.mux8 port map(mux_input_247, sel_mux, data_out(247));
inst_mux_248: entity work.mux8 port map(mux_input_248, sel_mux, data_out(248));
inst_mux_249: entity work.mux8 port map(mux_input_249, sel_mux, data_out(249));
inst_mux_250: entity work.mux8 port map(mux_input_250, sel_mux, data_out(250));
inst_mux_251: entity work.mux8 port map(mux_input_251, sel_mux, data_out(251));
inst_mux_252: entity work.mux8 port map(mux_input_252, sel_mux, data_out(252));
inst_mux_253: entity work.mux8 port map(mux_input_253, sel_mux, data_out(253));
inst_mux_254: entity work.mux8 port map(mux_input_254, sel_mux, data_out(254));
inst_mux_255: entity work.mux8 port map(mux_input_255, sel_mux, data_out(255));
end architecture;
