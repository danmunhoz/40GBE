------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 3.5
--  \   \         Application : 7 Series FPGAs Transceivers Wizard 
--  /   /         Filename : gtwizard_0_support.vhd
-- /___/   /\      
-- \   \  /  \ 
--  \___\/\___\
--
--  Description : This module instantiates the modules required for
--                reset and initialisation of the Transceiver
--
-- Module gtwizard_0_support
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;
--***********************************Entity Declaration************************

entity gtwizard_0_support is
generic
(
    EXAMPLE_SIM_GTRESET_SPEEDUP             : string    := "TRUE";     -- simulation setting for GT SecureIP model
    STABLE_CLOCK_PERIOD                     : integer   := 10  

);
port
(
    SOFT_RESET_TX_IN                        : in   std_logic;
    SOFT_RESET_RX_IN                        : in   std_logic;
    DONT_RESET_ON_DATA_ERROR_IN             : in   std_logic;
    Q8_CLK0_GTREFCLK_PAD_N_IN               : in   std_logic;
    Q8_CLK0_GTREFCLK_PAD_P_IN               : in   std_logic;
    Q8_CLK0_GTREFCLK_OUT                    : out  std_logic;
    GT0_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_DATA_VALID_IN                       : in   std_logic;
    GT0_TX_MMCM_LOCK_OUT                    : out  std_logic;
    GT0_RX_MMCM_LOCK_OUT                    : out  std_logic;
    GT1_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT1_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT1_DATA_VALID_IN                       : in   std_logic;
    GT1_TX_MMCM_LOCK_OUT                    : out  std_logic;
    GT1_RX_MMCM_LOCK_OUT                    : out  std_logic;
    GT2_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT2_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT2_DATA_VALID_IN                       : in   std_logic;
    GT2_TX_MMCM_LOCK_OUT                    : out  std_logic;
    GT2_RX_MMCM_LOCK_OUT                    : out  std_logic;
    GT3_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT3_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT3_DATA_VALID_IN                       : in   std_logic;
    GT3_TX_MMCM_LOCK_OUT                    : out  std_logic;
    GT3_RX_MMCM_LOCK_OUT                    : out  std_logic;
 
    GT0_TXUSRCLK_OUT                        : out  std_logic;
    GT0_TXUSRCLK2_OUT                       : out  std_logic;
    GT0_RXUSRCLK_OUT                        : out  std_logic;
    GT0_RXUSRCLK2_OUT                       : out  std_logic;
 
    GT1_TXUSRCLK_OUT                        : out  std_logic;
    GT1_TXUSRCLK2_OUT                       : out  std_logic;
    GT1_RXUSRCLK_OUT                        : out  std_logic;
    GT1_RXUSRCLK2_OUT                       : out  std_logic;
 
    GT2_TXUSRCLK_OUT                        : out  std_logic;
    GT2_TXUSRCLK2_OUT                       : out  std_logic;
    GT2_RXUSRCLK_OUT                        : out  std_logic;
    GT2_RXUSRCLK2_OUT                       : out  std_logic;
 
    GT3_TXUSRCLK_OUT                        : out  std_logic;
    GT3_TXUSRCLK2_OUT                       : out  std_logic;
    GT3_RXUSRCLK_OUT                        : out  std_logic;
    GT3_RXUSRCLK2_OUT                       : out  std_logic;

    --_________________________________________________________________________
    --GT0  (X1Y36)
    --____________________________CHANNEL PORTS________________________________
    ------------------------------- Loopback Ports -----------------------------
    gt0_loopback_in                         : in   std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt0_eyescanreset_in                     : in   std_logic;
    gt0_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt0_eyescandataerror_out                : out  std_logic;
    gt0_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt0_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt0_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------- Receive Ports - Pattern Checker Ports ------------------
    gt0_rxprbserr_out                       : out  std_logic;
    gt0_rxprbssel_in                        : in   std_logic_vector(2 downto 0);
    ------------------- Receive Ports - Pattern Checker ports ------------------
    gt0_rxprbscntreset_in                   : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt0_gthrxn_in                           : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt0_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt0_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    ---------------------- Receive Ports - RX Gearbox Ports --------------------
    gt0_rxdatavalid_out                     : out  std_logic;
    gt0_rxheader_out                        : out  std_logic_vector(1 downto 0);
    gt0_rxheadervalid_out                   : out  std_logic;
    --------------------- Receive Ports - RX Gearbox Ports  --------------------
    gt0_rxgearboxslip_in                    : in   std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt0_gtrxreset_in                        : in   std_logic;
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt0_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt0_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt0_gttxreset_in                        : in   std_logic;
    gt0_txuserrdy_in                        : in   std_logic;
    -------------- Transmit Ports - 64b66b and 64b67b Gearbox Ports ------------
    gt0_txheader_in                         : in   std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - Pattern Generator Ports ----------------
    gt0_txprbsforceerr_in                   : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt0_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt0_gthtxn_out                          : out  std_logic;
    gt0_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt0_txoutclkfabric_out                  : out  std_logic;
    gt0_txoutclkpcs_out                     : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    gt0_txsequence_in                       : in   std_logic_vector(6 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt0_txresetdone_out                     : out  std_logic;
    ------------------ Transmit Ports - pattern Generator Ports ----------------
    gt0_txprbssel_in                        : in   std_logic_vector(2 downto 0);

    --GT1  (X1Y37)
    --____________________________CHANNEL PORTS________________________________
    ------------------------------- Loopback Ports -----------------------------
    gt1_loopback_in                         : in   std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt1_eyescanreset_in                     : in   std_logic;
    gt1_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt1_eyescandataerror_out                : out  std_logic;
    gt1_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt1_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt1_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------- Receive Ports - Pattern Checker Ports ------------------
    gt1_rxprbserr_out                       : out  std_logic;
    gt1_rxprbssel_in                        : in   std_logic_vector(2 downto 0);
    ------------------- Receive Ports - Pattern Checker ports ------------------
    gt1_rxprbscntreset_in                   : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt1_gthrxn_in                           : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt1_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt1_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    ---------------------- Receive Ports - RX Gearbox Ports --------------------
    gt1_rxdatavalid_out                     : out  std_logic;
    gt1_rxheader_out                        : out  std_logic_vector(1 downto 0);
    gt1_rxheadervalid_out                   : out  std_logic;
    --------------------- Receive Ports - RX Gearbox Ports  --------------------
    gt1_rxgearboxslip_in                    : in   std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt1_gtrxreset_in                        : in   std_logic;
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt1_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt1_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt1_gttxreset_in                        : in   std_logic;
    gt1_txuserrdy_in                        : in   std_logic;
    -------------- Transmit Ports - 64b66b and 64b67b Gearbox Ports ------------
    gt1_txheader_in                         : in   std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - Pattern Generator Ports ----------------
    gt1_txprbsforceerr_in                   : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt1_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt1_gthtxn_out                          : out  std_logic;
    gt1_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt1_txoutclkfabric_out                  : out  std_logic;
    gt1_txoutclkpcs_out                     : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    gt1_txsequence_in                       : in   std_logic_vector(6 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt1_txresetdone_out                     : out  std_logic;
    ------------------ Transmit Ports - pattern Generator Ports ----------------
    gt1_txprbssel_in                        : in   std_logic_vector(2 downto 0);

    --GT2  (X1Y38)
    --____________________________CHANNEL PORTS________________________________
    ------------------------------- Loopback Ports -----------------------------
    gt2_loopback_in                         : in   std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt2_eyescanreset_in                     : in   std_logic;
    gt2_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt2_eyescandataerror_out                : out  std_logic;
    gt2_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt2_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt2_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------- Receive Ports - Pattern Checker Ports ------------------
    gt2_rxprbserr_out                       : out  std_logic;
    gt2_rxprbssel_in                        : in   std_logic_vector(2 downto 0);
    ------------------- Receive Ports - Pattern Checker ports ------------------
    gt2_rxprbscntreset_in                   : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt2_gthrxn_in                           : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt2_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt2_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    ---------------------- Receive Ports - RX Gearbox Ports --------------------
    gt2_rxdatavalid_out                     : out  std_logic;
    gt2_rxheader_out                        : out  std_logic_vector(1 downto 0);
    gt2_rxheadervalid_out                   : out  std_logic;
    --------------------- Receive Ports - RX Gearbox Ports  --------------------
    gt2_rxgearboxslip_in                    : in   std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt2_gtrxreset_in                        : in   std_logic;
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt2_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt2_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt2_gttxreset_in                        : in   std_logic;
    gt2_txuserrdy_in                        : in   std_logic;
    -------------- Transmit Ports - 64b66b and 64b67b Gearbox Ports ------------
    gt2_txheader_in                         : in   std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - Pattern Generator Ports ----------------
    gt2_txprbsforceerr_in                   : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt2_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt2_gthtxn_out                          : out  std_logic;
    gt2_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt2_txoutclkfabric_out                  : out  std_logic;
    gt2_txoutclkpcs_out                     : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    gt2_txsequence_in                       : in   std_logic_vector(6 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt2_txresetdone_out                     : out  std_logic;
    ------------------ Transmit Ports - pattern Generator Ports ----------------
    gt2_txprbssel_in                        : in   std_logic_vector(2 downto 0);

    --GT3  (X1Y39)
    --____________________________CHANNEL PORTS________________________________
    ------------------------------- Loopback Ports -----------------------------
    gt3_loopback_in                         : in   std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt3_eyescanreset_in                     : in   std_logic;
    gt3_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt3_eyescandataerror_out                : out  std_logic;
    gt3_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt3_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt3_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------- Receive Ports - Pattern Checker Ports ------------------
    gt3_rxprbserr_out                       : out  std_logic;
    gt3_rxprbssel_in                        : in   std_logic_vector(2 downto 0);
    ------------------- Receive Ports - Pattern Checker ports ------------------
    gt3_rxprbscntreset_in                   : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt3_gthrxn_in                           : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt3_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt3_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    ---------------------- Receive Ports - RX Gearbox Ports --------------------
    gt3_rxdatavalid_out                     : out  std_logic;
    gt3_rxheader_out                        : out  std_logic_vector(1 downto 0);
    gt3_rxheadervalid_out                   : out  std_logic;
    --------------------- Receive Ports - RX Gearbox Ports  --------------------
    gt3_rxgearboxslip_in                    : in   std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt3_gtrxreset_in                        : in   std_logic;
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt3_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt3_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt3_gttxreset_in                        : in   std_logic;
    gt3_txuserrdy_in                        : in   std_logic;
    -------------- Transmit Ports - 64b66b and 64b67b Gearbox Ports ------------
    gt3_txheader_in                         : in   std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - Pattern Generator Ports ----------------
    gt3_txprbsforceerr_in                   : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt3_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt3_gthtxn_out                          : out  std_logic;
    gt3_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt3_txoutclkfabric_out                  : out  std_logic;
    gt3_txoutclkpcs_out                     : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    gt3_txsequence_in                       : in   std_logic_vector(6 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt3_txresetdone_out                     : out  std_logic;
    ------------------ Transmit Ports - pattern Generator Ports ----------------
    gt3_txprbssel_in                        : in   std_logic_vector(2 downto 0);

    --____________________________COMMON PORTS________________________________
    GT0_QPLLLOCK_OUT : out std_logic;
    GT0_QPLLREFCLKLOST_OUT  : out std_logic;
    GT0_QPLLOUTCLK_OUT  : out std_logic;
    GT0_QPLLOUTREFCLK_OUT : out std_logic;
    
 
    

    sysclk_in        : in std_logic

);

end gtwizard_0_support;
    
architecture RTL of gtwizard_0_support is
attribute DowngradeIPIdentifiedWarnings: string;
attribute DowngradeIPIdentifiedWarnings of RTL : architecture is "yes";

--**************************Component Declarations*****************************

component gtwizard_0
 
port
(
    SYSCLK_IN                               : in   std_logic;
    SOFT_RESET_TX_IN                        : in   std_logic;
    SOFT_RESET_RX_IN                        : in   std_logic;
    DONT_RESET_ON_DATA_ERROR_IN             : in   std_logic;
    GT0_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_DATA_VALID_IN                       : in   std_logic;
    GT0_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT0_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT0_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT0_RX_MMCM_RESET_OUT                   : out  std_logic;
    GT1_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT1_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT1_DATA_VALID_IN                       : in   std_logic;
    GT1_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT1_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT1_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT1_RX_MMCM_RESET_OUT                   : out  std_logic;
    GT2_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT2_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT2_DATA_VALID_IN                       : in   std_logic;
    GT2_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT2_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT2_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT2_RX_MMCM_RESET_OUT                   : out  std_logic;
    GT3_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT3_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT3_DATA_VALID_IN                       : in   std_logic;
    GT3_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT3_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT3_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT3_RX_MMCM_RESET_OUT                   : out  std_logic;

    --_________________________________________________________________________
    --GT0  (X1Y36)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt0_drpclk_in                           : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    gt0_loopback_in                         : in   std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt0_eyescanreset_in                     : in   std_logic;
    gt0_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt0_eyescandataerror_out                : out  std_logic;
    gt0_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt0_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt0_rxusrclk_in                         : in   std_logic;
    gt0_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt0_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------- Receive Ports - Pattern Checker Ports ------------------
    gt0_rxprbserr_out                       : out  std_logic;
    gt0_rxprbssel_in                        : in   std_logic_vector(2 downto 0);
    ------------------- Receive Ports - Pattern Checker ports ------------------
    gt0_rxprbscntreset_in                   : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt0_gthrxn_in                           : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt0_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt0_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt0_rxoutclk_out                        : out  std_logic;
    ---------------------- Receive Ports - RX Gearbox Ports --------------------
    gt0_rxdatavalid_out                     : out  std_logic;
    gt0_rxheader_out                        : out  std_logic_vector(1 downto 0);
    gt0_rxheadervalid_out                   : out  std_logic;
    --------------------- Receive Ports - RX Gearbox Ports  --------------------
    gt0_rxgearboxslip_in                    : in   std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt0_gtrxreset_in                        : in   std_logic;
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt0_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt0_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt0_gttxreset_in                        : in   std_logic;
    gt0_txuserrdy_in                        : in   std_logic;
    -------------- Transmit Ports - 64b66b and 64b67b Gearbox Ports ------------
    gt0_txheader_in                         : in   std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt0_txusrclk_in                         : in   std_logic;
    gt0_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - Pattern Generator Ports ----------------
    gt0_txprbsforceerr_in                   : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt0_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt0_gthtxn_out                          : out  std_logic;
    gt0_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt0_txoutclk_out                        : out  std_logic;
    gt0_txoutclkfabric_out                  : out  std_logic;
    gt0_txoutclkpcs_out                     : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    gt0_txsequence_in                       : in   std_logic_vector(6 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt0_txresetdone_out                     : out  std_logic;
    ------------------ Transmit Ports - pattern Generator Ports ----------------
    gt0_txprbssel_in                        : in   std_logic_vector(2 downto 0);

    --GT1  (X1Y37)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt1_drpclk_in                           : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    gt1_loopback_in                         : in   std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt1_eyescanreset_in                     : in   std_logic;
    gt1_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt1_eyescandataerror_out                : out  std_logic;
    gt1_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt1_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt1_rxusrclk_in                         : in   std_logic;
    gt1_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt1_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------- Receive Ports - Pattern Checker Ports ------------------
    gt1_rxprbserr_out                       : out  std_logic;
    gt1_rxprbssel_in                        : in   std_logic_vector(2 downto 0);
    ------------------- Receive Ports - Pattern Checker ports ------------------
    gt1_rxprbscntreset_in                   : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt1_gthrxn_in                           : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt1_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt1_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt1_rxoutclk_out                        : out  std_logic;
    ---------------------- Receive Ports - RX Gearbox Ports --------------------
    gt1_rxdatavalid_out                     : out  std_logic;
    gt1_rxheader_out                        : out  std_logic_vector(1 downto 0);
    gt1_rxheadervalid_out                   : out  std_logic;
    --------------------- Receive Ports - RX Gearbox Ports  --------------------
    gt1_rxgearboxslip_in                    : in   std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt1_gtrxreset_in                        : in   std_logic;
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt1_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt1_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt1_gttxreset_in                        : in   std_logic;
    gt1_txuserrdy_in                        : in   std_logic;
    -------------- Transmit Ports - 64b66b and 64b67b Gearbox Ports ------------
    gt1_txheader_in                         : in   std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt1_txusrclk_in                         : in   std_logic;
    gt1_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - Pattern Generator Ports ----------------
    gt1_txprbsforceerr_in                   : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt1_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt1_gthtxn_out                          : out  std_logic;
    gt1_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt1_txoutclk_out                        : out  std_logic;
    gt1_txoutclkfabric_out                  : out  std_logic;
    gt1_txoutclkpcs_out                     : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    gt1_txsequence_in                       : in   std_logic_vector(6 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt1_txresetdone_out                     : out  std_logic;
    ------------------ Transmit Ports - pattern Generator Ports ----------------
    gt1_txprbssel_in                        : in   std_logic_vector(2 downto 0);

    --GT2  (X1Y38)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt2_drpclk_in                           : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    gt2_loopback_in                         : in   std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt2_eyescanreset_in                     : in   std_logic;
    gt2_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt2_eyescandataerror_out                : out  std_logic;
    gt2_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt2_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt2_rxusrclk_in                         : in   std_logic;
    gt2_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt2_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------- Receive Ports - Pattern Checker Ports ------------------
    gt2_rxprbserr_out                       : out  std_logic;
    gt2_rxprbssel_in                        : in   std_logic_vector(2 downto 0);
    ------------------- Receive Ports - Pattern Checker ports ------------------
    gt2_rxprbscntreset_in                   : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt2_gthrxn_in                           : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt2_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt2_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt2_rxoutclk_out                        : out  std_logic;
    ---------------------- Receive Ports - RX Gearbox Ports --------------------
    gt2_rxdatavalid_out                     : out  std_logic;
    gt2_rxheader_out                        : out  std_logic_vector(1 downto 0);
    gt2_rxheadervalid_out                   : out  std_logic;
    --------------------- Receive Ports - RX Gearbox Ports  --------------------
    gt2_rxgearboxslip_in                    : in   std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt2_gtrxreset_in                        : in   std_logic;
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt2_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt2_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt2_gttxreset_in                        : in   std_logic;
    gt2_txuserrdy_in                        : in   std_logic;
    -------------- Transmit Ports - 64b66b and 64b67b Gearbox Ports ------------
    gt2_txheader_in                         : in   std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt2_txusrclk_in                         : in   std_logic;
    gt2_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - Pattern Generator Ports ----------------
    gt2_txprbsforceerr_in                   : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt2_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt2_gthtxn_out                          : out  std_logic;
    gt2_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt2_txoutclk_out                        : out  std_logic;
    gt2_txoutclkfabric_out                  : out  std_logic;
    gt2_txoutclkpcs_out                     : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    gt2_txsequence_in                       : in   std_logic_vector(6 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt2_txresetdone_out                     : out  std_logic;
    ------------------ Transmit Ports - pattern Generator Ports ----------------
    gt2_txprbssel_in                        : in   std_logic_vector(2 downto 0);

    --GT3  (X1Y39)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt3_drpclk_in                           : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    gt3_loopback_in                         : in   std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    gt3_eyescanreset_in                     : in   std_logic;
    gt3_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt3_eyescandataerror_out                : out  std_logic;
    gt3_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt3_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt3_rxusrclk_in                         : in   std_logic;
    gt3_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt3_rxdata_out                          : out  std_logic_vector(63 downto 0);
    ------------------- Receive Ports - Pattern Checker Ports ------------------
    gt3_rxprbserr_out                       : out  std_logic;
    gt3_rxprbssel_in                        : in   std_logic_vector(2 downto 0);
    ------------------- Receive Ports - Pattern Checker ports ------------------
    gt3_rxprbscntreset_in                   : in   std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt3_gthrxn_in                           : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt3_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt3_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt3_rxoutclk_out                        : out  std_logic;
    ---------------------- Receive Ports - RX Gearbox Ports --------------------
    gt3_rxdatavalid_out                     : out  std_logic;
    gt3_rxheader_out                        : out  std_logic_vector(1 downto 0);
    gt3_rxheadervalid_out                   : out  std_logic;
    --------------------- Receive Ports - RX Gearbox Ports  --------------------
    gt3_rxgearboxslip_in                    : in   std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt3_gtrxreset_in                        : in   std_logic;
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt3_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt3_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt3_gttxreset_in                        : in   std_logic;
    gt3_txuserrdy_in                        : in   std_logic;
    -------------- Transmit Ports - 64b66b and 64b67b Gearbox Ports ------------
    gt3_txheader_in                         : in   std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt3_txusrclk_in                         : in   std_logic;
    gt3_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - Pattern Generator Ports ----------------
    gt3_txprbsforceerr_in                   : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt3_txdata_in                           : in   std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt3_gthtxn_out                          : out  std_logic;
    gt3_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt3_txoutclk_out                        : out  std_logic;
    gt3_txoutclkfabric_out                  : out  std_logic;
    gt3_txoutclkpcs_out                     : out  std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    gt3_txsequence_in                       : in   std_logic_vector(6 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt3_txresetdone_out                     : out  std_logic;
    ------------------ Transmit Ports - pattern Generator Ports ----------------
    gt3_txprbssel_in                        : in   std_logic_vector(2 downto 0);


    --____________________________COMMON PORTS________________________________
    GT0_QPLLLOCK_IN : in std_logic;
    GT0_QPLLREFCLKLOST_IN  : in std_logic;
    GT0_QPLLRESET_OUT  : out std_logic;
    GT0_QPLLOUTCLK_IN  : in std_logic;
    GT0_QPLLOUTREFCLK_IN : in std_logic 

);

end component;

component gtwizard_0_common_reset  
generic
(
      STABLE_CLOCK_PERIOD      : integer := 8        -- Period of the stable clock driving this state-machine, unit is [ns]
   );
port
   (    
      STABLE_CLOCK             : in std_logic;             --Stable Clock, either a stable clock from the PCB
      SOFT_RESET               : in std_logic;               --User Reset, can be pulled any time
      COMMON_RESET             : out std_logic  --Reset QPLL
   );
end component;

component gtwizard_0_common 
generic
(
    -- Simulation attributes
    WRAPPER_SIM_GTRESET_SPEEDUP     : string     :=  "FALSE" ;       -- Set to "TRUE" to speed up sim reset
    SIM_QPLLREFCLK_SEL              :bit_vector  := "001"
 
);
port
(
    QPLLREFCLKSEL_IN   : in std_logic_vector(2 downto 0);
    GTREFCLK0_IN : in std_logic;
    GTREFCLK1_IN      : in std_logic;
    QPLLLOCK_OUT : out std_logic;
    QPLLLOCKDETCLK_IN : in std_logic;
    QPLLOUTCLK_OUT : out std_logic;
    QPLLOUTREFCLK_OUT : out std_logic;
    QPLLREFCLKLOST_OUT : out std_logic;    
    QPLLRESET_IN : in std_logic

);

end component;
component gtwizard_0_GT_USRCLK_SOURCE 
port
(
 
    GT0_TXUSRCLK_OUT             : out std_logic;
    GT0_TXUSRCLK2_OUT            : out std_logic;
    GT0_TXOUTCLK_IN              : in  std_logic;
    GT0_TXCLK_LOCK_OUT           : out std_logic;
    GT0_TX_MMCM_RESET_IN         : in std_logic;
    GT0_RXUSRCLK_OUT             : out std_logic;
    GT0_RXUSRCLK2_OUT            : out std_logic;
    GT0_RXOUTCLK_IN              : in  std_logic;
    GT0_RXCLK_LOCK_OUT           : out std_logic;
    GT0_RX_MMCM_RESET_IN         : in std_logic;
 
    GT1_TXUSRCLK_OUT             : out std_logic;
    GT1_TXUSRCLK2_OUT            : out std_logic;
    GT1_TXOUTCLK_IN              : in  std_logic;
    GT1_TXCLK_LOCK_OUT           : out std_logic;
    GT1_TX_MMCM_RESET_IN         : in std_logic;
    GT1_RXUSRCLK_OUT             : out std_logic;
    GT1_RXUSRCLK2_OUT            : out std_logic;
    GT1_RXOUTCLK_IN              : in  std_logic;
    GT1_RXCLK_LOCK_OUT           : out std_logic;
    GT1_RX_MMCM_RESET_IN         : in std_logic;
 
    GT2_TXUSRCLK_OUT             : out std_logic;
    GT2_TXUSRCLK2_OUT            : out std_logic;
    GT2_TXOUTCLK_IN              : in  std_logic;
    GT2_TXCLK_LOCK_OUT           : out std_logic;
    GT2_TX_MMCM_RESET_IN         : in std_logic;
    GT2_RXUSRCLK_OUT             : out std_logic;
    GT2_RXUSRCLK2_OUT            : out std_logic;
    GT2_RXOUTCLK_IN              : in  std_logic;
    GT2_RXCLK_LOCK_OUT           : out std_logic;
    GT2_RX_MMCM_RESET_IN         : in std_logic;
 
    GT3_TXUSRCLK_OUT             : out std_logic;
    GT3_TXUSRCLK2_OUT            : out std_logic;
    GT3_TXOUTCLK_IN              : in  std_logic;
    GT3_TXCLK_LOCK_OUT           : out std_logic;
    GT3_TX_MMCM_RESET_IN         : in std_logic;
    GT3_RXUSRCLK_OUT             : out std_logic;
    GT3_RXUSRCLK2_OUT            : out std_logic;
    GT3_RXOUTCLK_IN              : in  std_logic;
    GT3_RXCLK_LOCK_OUT           : out std_logic;
    GT3_RX_MMCM_RESET_IN         : in std_logic;
    Q8_CLK0_GTREFCLK_PAD_N_IN               : in   std_logic;
    Q8_CLK0_GTREFCLK_PAD_P_IN               : in   std_logic;
    Q8_CLK0_GTREFCLK_OUT                    : out  std_logic
);
end component;

--***********************************Parameter Declarations********************

    constant DLY : time := 1 ns;

--************************** Register Declarations ****************************

    signal   gt0_txfsmresetdone_i            : std_logic;
signal   gt0_rxfsmresetdone_i            : std_logic;
    signal   gt0_txfsmresetdone_r            : std_logic;
    signal   gt0_txfsmresetdone_r2           : std_logic;
signal   gt0_rxresetdone_r               : std_logic;
signal   gt0_rxresetdone_r2              : std_logic;
signal   gt0_rxresetdone_r3              : std_logic;

--***************************** Register Declarations *****************************
    signal   gt0_txseq_counter_r      :   unsigned(8 downto 0);
signal   gt0_txheader_r           :   std_logic_vector(1 downto 0);
signal   gt0_extend_reset_r       :   std_logic_vector(3 downto 0);
signal   gt0_pause_data_valid_r   :   std_logic;

    signal   gt1_txfsmresetdone_i            : std_logic;
signal   gt1_rxfsmresetdone_i            : std_logic;
    signal   gt1_txfsmresetdone_r            : std_logic;
    signal   gt1_txfsmresetdone_r2           : std_logic;
signal   gt1_rxresetdone_r               : std_logic;
signal   gt1_rxresetdone_r2              : std_logic;
signal   gt1_rxresetdone_r3              : std_logic;

--***************************** Register Declarations *****************************
    signal   gt1_txseq_counter_r      :   unsigned(8 downto 0);
signal   gt1_txheader_r           :   std_logic_vector(1 downto 0);
signal   gt1_extend_reset_r       :   std_logic_vector(3 downto 0);
signal   gt1_pause_data_valid_r   :   std_logic;

    signal   gt2_txfsmresetdone_i            : std_logic;
signal   gt2_rxfsmresetdone_i            : std_logic;
    signal   gt2_txfsmresetdone_r            : std_logic;
    signal   gt2_txfsmresetdone_r2           : std_logic;
signal   gt2_rxresetdone_r               : std_logic;
signal   gt2_rxresetdone_r2              : std_logic;
signal   gt2_rxresetdone_r3              : std_logic;

--***************************** Register Declarations *****************************
    signal   gt2_txseq_counter_r      :   unsigned(8 downto 0);
signal   gt2_txheader_r           :   std_logic_vector(1 downto 0);
signal   gt2_extend_reset_r       :   std_logic_vector(3 downto 0);
signal   gt2_pause_data_valid_r   :   std_logic;

    signal   gt3_txfsmresetdone_i            : std_logic;
signal   gt3_rxfsmresetdone_i            : std_logic;
    signal   gt3_txfsmresetdone_r            : std_logic;
    signal   gt3_txfsmresetdone_r2           : std_logic;
signal   gt3_rxresetdone_r               : std_logic;
signal   gt3_rxresetdone_r2              : std_logic;
signal   gt3_rxresetdone_r3              : std_logic;

--***************************** Register Declarations *****************************
    signal   gt3_txseq_counter_r      :   unsigned(8 downto 0);
signal   gt3_txheader_r           :   std_logic_vector(1 downto 0);
signal   gt3_extend_reset_r       :   std_logic_vector(3 downto 0);
signal   gt3_pause_data_valid_r   :   std_logic;

signal   reset_pulse                     : std_logic_vector(3 downto 0);
    signal   reset_counter  :   unsigned(5 downto 0) := "000000";


--**************************** Wire Declarations ******************************
    -------------------------- GT Wrapper Wires ------------------------------
    --________________________________________________________________________
    --________________________________________________________________________
    --GT0  (X1Y36)

    ------------------------------- Loopback Ports -----------------------------
    signal  gt0_loopback_i                  : std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt0_eyescanreset_i              : std_logic;
    signal  gt0_rxuserrdy_i                 : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt0_eyescandataerror_i          : std_logic;
    signal  gt0_eyescantrigger_i            : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt0_dmonitorout_i               : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt0_rxdata_i                    : std_logic_vector(63 downto 0);
    ------------------- Receive Ports - Pattern Checker Ports ------------------
    signal  gt0_rxprbserr_i                 : std_logic;
    signal  gt0_rxprbssel_i                 : std_logic_vector(2 downto 0);
    ------------------- Receive Ports - Pattern Checker ports ------------------
    signal  gt0_rxprbscntreset_i            : std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt0_gthrxn_i                    : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt0_rxdfeagchold_i              : std_logic;
    signal  gt0_rxdfelfhold_i               : std_logic;
    signal  gt0_rxmonitorout_i              : std_logic_vector(6 downto 0);
    signal  gt0_rxmonitorsel_i              : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt0_rxoutclk_i                  : std_logic;
    ---------------------- Receive Ports - RX Gearbox Ports --------------------
    signal  gt0_rxdatavalid_i               : std_logic;
    signal  gt0_rxheader_i                  : std_logic_vector(1 downto 0);
    signal  gt0_rxheadervalid_i             : std_logic;
    --------------------- Receive Ports - RX Gearbox Ports  --------------------
    signal  gt0_rxgearboxslip_i             : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt0_gtrxreset_i                 : std_logic;
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt0_gthrxp_i                    : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt0_rxresetdone_i               : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt0_gttxreset_i                 : std_logic;
    signal  gt0_txuserrdy_i                 : std_logic;
    -------------- Transmit Ports - 64b66b and 64b67b Gearbox Ports ------------
    signal  gt0_txheader_i                  : std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - Pattern Generator Ports ----------------
    signal  gt0_txprbsforceerr_i            : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt0_txdata_i                    : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt0_gthtxn_i                    : std_logic;
    signal  gt0_gthtxp_i                    : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt0_txoutclk_i                  : std_logic;
    signal  gt0_txoutclkfabric_i            : std_logic;
    signal  gt0_txoutclkpcs_i               : std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    signal  gt0_txsequence_i                : std_logic_vector(6 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt0_txresetdone_i               : std_logic;
    ------------------ Transmit Ports - pattern Generator Ports ----------------
    signal  gt0_txprbssel_i                 : std_logic_vector(2 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT1  (X1Y37)

    ------------------------------- Loopback Ports -----------------------------
    signal  gt1_loopback_i                  : std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt1_eyescanreset_i              : std_logic;
    signal  gt1_rxuserrdy_i                 : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt1_eyescandataerror_i          : std_logic;
    signal  gt1_eyescantrigger_i            : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt1_dmonitorout_i               : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt1_rxdata_i                    : std_logic_vector(63 downto 0);
    ------------------- Receive Ports - Pattern Checker Ports ------------------
    signal  gt1_rxprbserr_i                 : std_logic;
    signal  gt1_rxprbssel_i                 : std_logic_vector(2 downto 0);
    ------------------- Receive Ports - Pattern Checker ports ------------------
    signal  gt1_rxprbscntreset_i            : std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt1_gthrxn_i                    : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt1_rxdfeagchold_i              : std_logic;
    signal  gt1_rxdfelfhold_i               : std_logic;
    signal  gt1_rxmonitorout_i              : std_logic_vector(6 downto 0);
    signal  gt1_rxmonitorsel_i              : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt1_rxoutclk_i                  : std_logic;
    ---------------------- Receive Ports - RX Gearbox Ports --------------------
    signal  gt1_rxdatavalid_i               : std_logic;
    signal  gt1_rxheader_i                  : std_logic_vector(1 downto 0);
    signal  gt1_rxheadervalid_i             : std_logic;
    --------------------- Receive Ports - RX Gearbox Ports  --------------------
    signal  gt1_rxgearboxslip_i             : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt1_gtrxreset_i                 : std_logic;
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt1_gthrxp_i                    : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt1_rxresetdone_i               : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt1_gttxreset_i                 : std_logic;
    signal  gt1_txuserrdy_i                 : std_logic;
    -------------- Transmit Ports - 64b66b and 64b67b Gearbox Ports ------------
    signal  gt1_txheader_i                  : std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - Pattern Generator Ports ----------------
    signal  gt1_txprbsforceerr_i            : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt1_txdata_i                    : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt1_gthtxn_i                    : std_logic;
    signal  gt1_gthtxp_i                    : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt1_txoutclk_i                  : std_logic;
    signal  gt1_txoutclkfabric_i            : std_logic;
    signal  gt1_txoutclkpcs_i               : std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    signal  gt1_txsequence_i                : std_logic_vector(6 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt1_txresetdone_i               : std_logic;
    ------------------ Transmit Ports - pattern Generator Ports ----------------
    signal  gt1_txprbssel_i                 : std_logic_vector(2 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT2  (X1Y38)

    ------------------------------- Loopback Ports -----------------------------
    signal  gt2_loopback_i                  : std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt2_eyescanreset_i              : std_logic;
    signal  gt2_rxuserrdy_i                 : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt2_eyescandataerror_i          : std_logic;
    signal  gt2_eyescantrigger_i            : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt2_dmonitorout_i               : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt2_rxdata_i                    : std_logic_vector(63 downto 0);
    ------------------- Receive Ports - Pattern Checker Ports ------------------
    signal  gt2_rxprbserr_i                 : std_logic;
    signal  gt2_rxprbssel_i                 : std_logic_vector(2 downto 0);
    ------------------- Receive Ports - Pattern Checker ports ------------------
    signal  gt2_rxprbscntreset_i            : std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt2_gthrxn_i                    : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt2_rxdfeagchold_i              : std_logic;
    signal  gt2_rxdfelfhold_i               : std_logic;
    signal  gt2_rxmonitorout_i              : std_logic_vector(6 downto 0);
    signal  gt2_rxmonitorsel_i              : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt2_rxoutclk_i                  : std_logic;
    ---------------------- Receive Ports - RX Gearbox Ports --------------------
    signal  gt2_rxdatavalid_i               : std_logic;
    signal  gt2_rxheader_i                  : std_logic_vector(1 downto 0);
    signal  gt2_rxheadervalid_i             : std_logic;
    --------------------- Receive Ports - RX Gearbox Ports  --------------------
    signal  gt2_rxgearboxslip_i             : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt2_gtrxreset_i                 : std_logic;
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt2_gthrxp_i                    : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt2_rxresetdone_i               : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt2_gttxreset_i                 : std_logic;
    signal  gt2_txuserrdy_i                 : std_logic;
    -------------- Transmit Ports - 64b66b and 64b67b Gearbox Ports ------------
    signal  gt2_txheader_i                  : std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - Pattern Generator Ports ----------------
    signal  gt2_txprbsforceerr_i            : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt2_txdata_i                    : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt2_gthtxn_i                    : std_logic;
    signal  gt2_gthtxp_i                    : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt2_txoutclk_i                  : std_logic;
    signal  gt2_txoutclkfabric_i            : std_logic;
    signal  gt2_txoutclkpcs_i               : std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    signal  gt2_txsequence_i                : std_logic_vector(6 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt2_txresetdone_i               : std_logic;
    ------------------ Transmit Ports - pattern Generator Ports ----------------
    signal  gt2_txprbssel_i                 : std_logic_vector(2 downto 0);

    --________________________________________________________________________
    --________________________________________________________________________
    --GT3  (X1Y39)

    ------------------------------- Loopback Ports -----------------------------
    signal  gt3_loopback_i                  : std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt3_eyescanreset_i              : std_logic;
    signal  gt3_rxuserrdy_i                 : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt3_eyescandataerror_i          : std_logic;
    signal  gt3_eyescantrigger_i            : std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    signal  gt3_dmonitorout_i               : std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt3_rxdata_i                    : std_logic_vector(63 downto 0);
    ------------------- Receive Ports - Pattern Checker Ports ------------------
    signal  gt3_rxprbserr_i                 : std_logic;
    signal  gt3_rxprbssel_i                 : std_logic_vector(2 downto 0);
    ------------------- Receive Ports - Pattern Checker ports ------------------
    signal  gt3_rxprbscntreset_i            : std_logic;
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt3_gthrxn_i                    : std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    signal  gt3_rxdfeagchold_i              : std_logic;
    signal  gt3_rxdfelfhold_i               : std_logic;
    signal  gt3_rxmonitorout_i              : std_logic_vector(6 downto 0);
    signal  gt3_rxmonitorsel_i              : std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt3_rxoutclk_i                  : std_logic;
    ---------------------- Receive Ports - RX Gearbox Ports --------------------
    signal  gt3_rxdatavalid_i               : std_logic;
    signal  gt3_rxheader_i                  : std_logic_vector(1 downto 0);
    signal  gt3_rxheadervalid_i             : std_logic;
    --------------------- Receive Ports - RX Gearbox Ports  --------------------
    signal  gt3_rxgearboxslip_i             : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt3_gtrxreset_i                 : std_logic;
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt3_gthrxp_i                    : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt3_rxresetdone_i               : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt3_gttxreset_i                 : std_logic;
    signal  gt3_txuserrdy_i                 : std_logic;
    -------------- Transmit Ports - 64b66b and 64b67b Gearbox Ports ------------
    signal  gt3_txheader_i                  : std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - Pattern Generator Ports ----------------
    signal  gt3_txprbsforceerr_i            : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt3_txdata_i                    : std_logic_vector(63 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt3_gthtxn_i                    : std_logic;
    signal  gt3_gthtxp_i                    : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt3_txoutclk_i                  : std_logic;
    signal  gt3_txoutclkfabric_i            : std_logic;
    signal  gt3_txoutclkpcs_i               : std_logic;
    --------------------- Transmit Ports - TX Gearbox Ports --------------------
    signal  gt3_txsequence_i                : std_logic_vector(6 downto 0);
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt3_txresetdone_i               : std_logic;
    ------------------ Transmit Ports - pattern Generator Ports ----------------
    signal  gt3_txprbssel_i                 : std_logic_vector(2 downto 0);

    --____________________________COMMON PORTS________________________________
    signal gt0_qplllock_i : std_logic;
    signal gt0_qpllrefclklost_i  : std_logic;
    signal gt0_qpllreset_i  : std_logic;
    signal gt0_qpllreset_t  : std_logic;
    signal gt0_qplloutclk_i  : std_logic;
    signal gt0_qplloutrefclk_i : std_logic;
  
    ------------------------------- Global Signals -----------------------------
    signal  gt0_tx_system_reset_c           : std_logic;
    signal  gt0_rx_system_reset_c           : std_logic;
    signal  gt1_tx_system_reset_c           : std_logic;
    signal  gt1_rx_system_reset_c           : std_logic;
    signal  gt2_tx_system_reset_c           : std_logic;
    signal  gt2_rx_system_reset_c           : std_logic;
    signal  gt3_tx_system_reset_c           : std_logic;
    signal  gt3_rx_system_reset_c           : std_logic;
    signal  tied_to_ground_i                : std_logic;
    signal  tied_to_ground_vec_i            : std_logic_vector(63 downto 0);
    signal  tied_to_vcc_i                   : std_logic;
    signal  tied_to_vcc_vec_i               : std_logic_vector(7 downto 0);
    signal  drpclk_in_i                     : std_logic;
    signal  sysclk_in_i                     : std_logic;
    signal   gt0_rx_reset_i           :   std_logic;
    signal   gt0_rx_reset_i1          :   std_logic;
    signal   gt0_rx_reset_i2          :   std_logic;
    signal   gt0_not_block_lock_i     :   std_logic;
    signal   gt0_scrambled_data_i     :   std_logic_vector(63 downto 0);
    signal   gt0_data_valid_i         :   std_logic;
    signal   gt0_data_valid_out_i     :   std_logic;
    signal   gt0_tx_reset_i           :   std_logic;
    signal   gt0_reset_r              :   std_logic;
    signal   gt1_rx_reset_i           :   std_logic;
    signal   gt1_rx_reset_i1          :   std_logic;
    signal   gt1_rx_reset_i2          :   std_logic;
    signal   gt1_not_block_lock_i     :   std_logic;
    signal   gt1_scrambled_data_i     :   std_logic_vector(63 downto 0);
    signal   gt1_data_valid_i         :   std_logic;
    signal   gt1_data_valid_out_i     :   std_logic;
    signal   gt1_tx_reset_i           :   std_logic;
    signal   gt1_reset_r              :   std_logic;
    signal   gt2_rx_reset_i           :   std_logic;
    signal   gt2_rx_reset_i1          :   std_logic;
    signal   gt2_rx_reset_i2          :   std_logic;
    signal   gt2_not_block_lock_i     :   std_logic;
    signal   gt2_scrambled_data_i     :   std_logic_vector(63 downto 0);
    signal   gt2_data_valid_i         :   std_logic;
    signal   gt2_data_valid_out_i     :   std_logic;
    signal   gt2_tx_reset_i           :   std_logic;
    signal   gt2_reset_r              :   std_logic;
    signal   gt3_rx_reset_i           :   std_logic;
    signal   gt3_rx_reset_i1          :   std_logic;
    signal   gt3_rx_reset_i2          :   std_logic;
    signal   gt3_not_block_lock_i     :   std_logic;
    signal   gt3_scrambled_data_i     :   std_logic_vector(63 downto 0);
    signal   gt3_data_valid_i         :   std_logic;
    signal   gt3_data_valid_out_i     :   std_logic;
    signal   gt3_tx_reset_i           :   std_logic;
    signal   gt3_reset_r              :   std_logic;
    signal  GTTXRESET_IN                    : std_logic;
    signal  GTRXRESET_IN                    : std_logic;
    signal  QPLLRESET_IN                    : std_logic;

    attribute keep: string;
   ------------------------------- User Clocks ---------------------------------
    signal    gt0_txusrclk_i                  : std_logic; 
    signal    gt0_txusrclk2_i                 : std_logic; 
    signal    gt0_rxusrclk_i                  : std_logic; 
    signal    gt0_rxusrclk2_i                 : std_logic; 
    
    
    
    
    signal    gt1_txusrclk_i                  : std_logic; 
    signal    gt1_txusrclk2_i                 : std_logic; 
    signal    gt1_rxusrclk_i                  : std_logic; 
    signal    gt1_rxusrclk2_i                 : std_logic; 
    
    
    
    
    signal    gt2_txusrclk_i                  : std_logic; 
    signal    gt2_txusrclk2_i                 : std_logic; 
    signal    gt2_rxusrclk_i                  : std_logic; 
    signal    gt2_rxusrclk2_i                 : std_logic; 
    
    
    
    
    signal    gt3_txusrclk_i                  : std_logic; 
    signal    gt3_txusrclk2_i                 : std_logic; 
    signal    gt3_rxusrclk_i                  : std_logic; 
    signal    gt3_rxusrclk2_i                 : std_logic; 
    
    
    
    
    signal    gt0_txmmcm_lock_i               : std_logic;
    signal    gt0_txmmcm_reset_i              : std_logic;
    signal    gt0_rxmmcm_lock_i               : std_logic; 
    signal    gt0_rxmmcm_reset_i              : std_logic;
    signal    gt1_txmmcm_lock_i               : std_logic;
    signal    gt1_txmmcm_reset_i              : std_logic;
    signal    gt1_rxmmcm_lock_i               : std_logic; 
    signal    gt1_rxmmcm_reset_i              : std_logic;
    signal    gt2_txmmcm_lock_i               : std_logic;
    signal    gt2_txmmcm_reset_i              : std_logic;
    signal    gt2_rxmmcm_lock_i               : std_logic; 
    signal    gt2_rxmmcm_reset_i              : std_logic;
    signal    gt3_txmmcm_lock_i               : std_logic;
    signal    gt3_txmmcm_reset_i              : std_logic;
    signal    gt3_rxmmcm_lock_i               : std_logic; 
    signal    gt3_rxmmcm_reset_i              : std_logic;
    ----------------------------- Reference Clocks ----------------------------
    
signal    q8_clk0_refclk_i                : std_logic;

signal commonreset_i : std_logic;
--**************************** Main Body of Code *******************************
begin

    --  Static signal Assigments
tied_to_ground_i                             <= '0';
tied_to_ground_vec_i                         <= x"0000000000000000";
tied_to_vcc_i                                <= '1';
tied_to_vcc_vec_i                            <= "11111111";

     GT0_TX_MMCM_LOCK_OUT <= gt0_txmmcm_lock_i;
    GT0_RX_MMCM_LOCK_OUT <= gt0_rxmmcm_lock_i;
     GT1_TX_MMCM_LOCK_OUT <= gt1_txmmcm_lock_i;
    GT1_RX_MMCM_LOCK_OUT <= gt1_rxmmcm_lock_i;
     GT2_TX_MMCM_LOCK_OUT <= gt2_txmmcm_lock_i;
    GT2_RX_MMCM_LOCK_OUT <= gt2_rxmmcm_lock_i;
     GT3_TX_MMCM_LOCK_OUT <= gt3_txmmcm_lock_i;
    GT3_RX_MMCM_LOCK_OUT <= gt3_rxmmcm_lock_i;
 
      gt0_qplllock_out  <= gt0_qplllock_i;
      gt0_qpllrefclklost_out <= gt0_qpllrefclklost_i;
     gt0_qpllreset_t <= commonreset_i or gt0_qpllreset_i;
     gt0_qplloutclk_out <= gt0_qplloutclk_i;
     gt0_qplloutrefclk_out <= gt0_qplloutrefclk_i;


 
      GT0_TXUSRCLK_OUT <= gt0_txusrclk_i; 
      GT0_TXUSRCLK2_OUT <= gt0_txusrclk2_i;
      GT0_RXUSRCLK_OUT <= gt0_rxusrclk_i;
      GT0_RXUSRCLK2_OUT <= gt0_rxusrclk2_i;
 
      GT1_TXUSRCLK_OUT <= gt1_txusrclk_i; 
      GT1_TXUSRCLK2_OUT <= gt1_txusrclk2_i;
      GT1_RXUSRCLK_OUT <= gt1_rxusrclk_i;
      GT1_RXUSRCLK2_OUT <= gt1_rxusrclk2_i;
 
      GT2_TXUSRCLK_OUT <= gt2_txusrclk_i; 
      GT2_TXUSRCLK2_OUT <= gt2_txusrclk2_i;
      GT2_RXUSRCLK_OUT <= gt2_rxusrclk_i;
      GT2_RXUSRCLK2_OUT <= gt2_rxusrclk2_i;
 
      GT3_TXUSRCLK_OUT <= gt3_txusrclk_i; 
      GT3_TXUSRCLK2_OUT <= gt3_txusrclk2_i;
      GT3_RXUSRCLK_OUT <= gt3_rxusrclk_i;
      GT3_RXUSRCLK2_OUT <= gt3_rxusrclk2_i;


    gt_usrclk_source : gtwizard_0_GT_USRCLK_SOURCE
    port map
   (
 
        GT0_TXUSRCLK_OUT                =>      gt0_txusrclk_i,
        GT0_TXUSRCLK2_OUT               =>      gt0_txusrclk2_i,
        GT0_TXOUTCLK_IN                 =>      gt0_txoutclk_i,
        GT0_TXCLK_LOCK_OUT              =>      gt0_txmmcm_lock_i,
        GT0_TX_MMCM_RESET_IN            =>      gt0_txmmcm_reset_i,
        GT0_RXUSRCLK_OUT                =>      gt0_rxusrclk_i,
        GT0_RXUSRCLK2_OUT               =>      gt0_rxusrclk2_i,
        GT0_RXOUTCLK_IN                 =>      gt0_rxoutclk_i,
        GT0_RXCLK_LOCK_OUT              =>      gt0_rxmmcm_lock_i,
        GT0_RX_MMCM_RESET_IN            =>      gt0_rxmmcm_reset_i,
 
        GT1_TXUSRCLK_OUT                =>      gt1_txusrclk_i,
        GT1_TXUSRCLK2_OUT               =>      gt1_txusrclk2_i,
        GT1_TXOUTCLK_IN                 =>      gt1_txoutclk_i,
        GT1_TXCLK_LOCK_OUT              =>      gt1_txmmcm_lock_i,
        GT1_TX_MMCM_RESET_IN            =>      gt1_txmmcm_reset_i,
        GT1_RXUSRCLK_OUT                =>      gt1_rxusrclk_i,
        GT1_RXUSRCLK2_OUT               =>      gt1_rxusrclk2_i,
        GT1_RXOUTCLK_IN                 =>      gt1_rxoutclk_i,
        GT1_RXCLK_LOCK_OUT              =>      gt1_rxmmcm_lock_i,
        GT1_RX_MMCM_RESET_IN            =>      gt1_rxmmcm_reset_i,
 
        GT2_TXUSRCLK_OUT                =>      gt2_txusrclk_i,
        GT2_TXUSRCLK2_OUT               =>      gt2_txusrclk2_i,
        GT2_TXOUTCLK_IN                 =>      gt2_txoutclk_i,
        GT2_TXCLK_LOCK_OUT              =>      gt2_txmmcm_lock_i,
        GT2_TX_MMCM_RESET_IN            =>      gt2_txmmcm_reset_i,
        GT2_RXUSRCLK_OUT                =>      gt2_rxusrclk_i,
        GT2_RXUSRCLK2_OUT               =>      gt2_rxusrclk2_i,
        GT2_RXOUTCLK_IN                 =>      gt2_rxoutclk_i,
        GT2_RXCLK_LOCK_OUT              =>      gt2_rxmmcm_lock_i,
        GT2_RX_MMCM_RESET_IN            =>      gt2_rxmmcm_reset_i,
 
        GT3_TXUSRCLK_OUT                =>      gt3_txusrclk_i,
        GT3_TXUSRCLK2_OUT               =>      gt3_txusrclk2_i,
        GT3_TXOUTCLK_IN                 =>      gt3_txoutclk_i,
        GT3_TXCLK_LOCK_OUT              =>      gt3_txmmcm_lock_i,
        GT3_TX_MMCM_RESET_IN            =>      gt3_txmmcm_reset_i,
        GT3_RXUSRCLK_OUT                =>      gt3_rxusrclk_i,
        GT3_RXUSRCLK2_OUT               =>      gt3_rxusrclk2_i,
        GT3_RXOUTCLK_IN                 =>      gt3_rxoutclk_i,
        GT3_RXCLK_LOCK_OUT              =>      gt3_rxmmcm_lock_i,
        GT3_RX_MMCM_RESET_IN            =>      gt3_rxmmcm_reset_i,
        Q8_CLK0_GTREFCLK_PAD_N_IN       =>      Q8_CLK0_GTREFCLK_PAD_N_IN,
        Q8_CLK0_GTREFCLK_PAD_P_IN       =>      Q8_CLK0_GTREFCLK_PAD_P_IN,
        Q8_CLK0_GTREFCLK_OUT            =>      q8_clk0_refclk_i

    );

    sysclk_in_i <= sysclk_in;
    Q8_CLK0_GTREFCLK_OUT <= q8_clk0_refclk_i;

    common0_i:gtwizard_0_common 
  generic map
  (
   WRAPPER_SIM_GTRESET_SPEEDUP => EXAMPLE_SIM_GTRESET_SPEEDUP,
   SIM_QPLLREFCLK_SEL => "001"
  )
 port map
   (
    QPLLREFCLKSEL_IN    => "001",
    GTREFCLK0_IN      => q8_clk0_refclk_i,
    GTREFCLK1_IN      => tied_to_ground_i,
    QPLLLOCK_OUT => gt0_qplllock_i,
    QPLLLOCKDETCLK_IN => sysclk_in_i,
    QPLLOUTCLK_OUT => gt0_qplloutclk_i,
    QPLLOUTREFCLK_OUT => gt0_qplloutrefclk_i,
    QPLLREFCLKLOST_OUT => gt0_qpllrefclklost_i,    
    QPLLRESET_IN => gt0_qpllreset_t

);

    common_reset_i:gtwizard_0_common_reset 
   generic map 
   (
      STABLE_CLOCK_PERIOD =>STABLE_CLOCK_PERIOD        -- Period of the stable clock driving this state-machine, unit is [ns]
   )
   port map
   (    
      STABLE_CLOCK => sysclk_in_i,             --Stable Clock, either a stable clock from the PCB
     
      SOFT_RESET => soft_reset_tx_in,               --User Reset, can be pulled any time
      COMMON_RESET => commonreset_i              --Reset QPLL
   );


    gtwizard_0_init_i : gtwizard_0
    port map
    (
        sysclk_in                       =>      sysclk_in_i,
        soft_reset_tx_in                =>      SOFT_RESET_TX_IN,
        soft_reset_rx_in                =>      SOFT_RESET_RX_IN,
        dont_reset_on_data_error_in     =>      DONT_RESET_ON_DATA_ERROR_IN,
        gt0_tx_mmcm_lock_in             =>      gt0_txmmcm_lock_i,
        gt0_tx_mmcm_reset_out           =>      gt0_txmmcm_reset_i,
        gt0_rx_mmcm_lock_in             =>      gt0_rxmmcm_lock_i,
        gt0_rx_mmcm_reset_out           =>      gt0_rxmmcm_reset_i,
        gt0_tx_fsm_reset_done_out       =>      gt0_tx_fsm_reset_done_out,
        gt0_rx_fsm_reset_done_out       =>      gt0_rx_fsm_reset_done_out,
        gt0_data_valid_in               =>      gt0_data_valid_in,
        gt1_tx_mmcm_lock_in             =>      gt1_txmmcm_lock_i,
        gt1_tx_mmcm_reset_out           =>      gt1_txmmcm_reset_i,
        gt1_rx_mmcm_lock_in             =>      gt1_rxmmcm_lock_i,
        gt1_rx_mmcm_reset_out           =>      gt1_rxmmcm_reset_i,
        gt1_tx_fsm_reset_done_out       =>      gt1_tx_fsm_reset_done_out,
        gt1_rx_fsm_reset_done_out       =>      gt1_rx_fsm_reset_done_out,
        gt1_data_valid_in               =>      gt1_data_valid_in,
        gt2_tx_mmcm_lock_in             =>      gt2_txmmcm_lock_i,
        gt2_tx_mmcm_reset_out           =>      gt2_txmmcm_reset_i,
        gt2_rx_mmcm_lock_in             =>      gt2_rxmmcm_lock_i,
        gt2_rx_mmcm_reset_out           =>      gt2_rxmmcm_reset_i,
        gt2_tx_fsm_reset_done_out       =>      gt2_tx_fsm_reset_done_out,
        gt2_rx_fsm_reset_done_out       =>      gt2_rx_fsm_reset_done_out,
        gt2_data_valid_in               =>      gt2_data_valid_in,
        gt3_tx_mmcm_lock_in             =>      gt3_txmmcm_lock_i,
        gt3_tx_mmcm_reset_out           =>      gt3_txmmcm_reset_i,
        gt3_rx_mmcm_lock_in             =>      gt3_rxmmcm_lock_i,
        gt3_rx_mmcm_reset_out           =>      gt3_rxmmcm_reset_i,
        gt3_tx_fsm_reset_done_out       =>      gt3_tx_fsm_reset_done_out,
        gt3_rx_fsm_reset_done_out       =>      gt3_rx_fsm_reset_done_out,
        gt3_data_valid_in               =>      gt3_data_valid_in,

        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT0  (X1Y36)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt0_drpclk_in                   =>      sysclk_in_i,
        ------------------------------- Loopback Ports -----------------------------
        gt0_loopback_in                 =>      gt0_loopback_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt0_eyescanreset_in             =>      gt0_eyescanreset_in,
        gt0_rxuserrdy_in                =>      gt0_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt0_eyescandataerror_out        =>      gt0_eyescandataerror_out,
        gt0_eyescantrigger_in           =>      gt0_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt0_dmonitorout_out             =>      gt0_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt0_rxusrclk_in                 =>      gt0_rxusrclk_i,
        gt0_rxusrclk2_in                =>      gt0_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt0_rxdata_out                  =>      gt0_rxdata_out,
        ------------------- Receive Ports - Pattern Checker Ports ------------------
        gt0_rxprbserr_out               =>      gt0_rxprbserr_out,
        gt0_rxprbssel_in                =>      gt0_rxprbssel_in,
        ------------------- Receive Ports - Pattern Checker ports ------------------
        gt0_rxprbscntreset_in           =>      gt0_rxprbscntreset_in,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt0_gthrxn_in                   =>      gt0_gthrxn_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt0_rxmonitorout_out            =>      gt0_rxmonitorout_out,
        gt0_rxmonitorsel_in             =>      gt0_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt0_rxoutclk_out                =>      gt0_rxoutclk_i,
        ---------------------- Receive Ports - RX Gearbox Ports --------------------
        gt0_rxdatavalid_out             =>      gt0_rxdatavalid_out,
        gt0_rxheader_out                =>      gt0_rxheader_out,
        gt0_rxheadervalid_out           =>      gt0_rxheadervalid_out,
        --------------------- Receive Ports - RX Gearbox Ports  --------------------
        gt0_rxgearboxslip_in            =>      gt0_rxgearboxslip_in,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt0_gtrxreset_in                =>      gt0_gtrxreset_in,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt0_gthrxp_in                   =>      gt0_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt0_rxresetdone_out             =>      gt0_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt0_gttxreset_in                =>      gt0_gttxreset_in,
        gt0_txuserrdy_in                =>      gt0_txuserrdy_in,
        -------------- Transmit Ports - 64b66b and 64b67b Gearbox Ports ------------
        gt0_txheader_in                 =>      gt0_txheader_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt0_txusrclk_in                 =>      gt0_txusrclk_i,
        gt0_txusrclk2_in                =>      gt0_txusrclk2_i,
        ------------------ Transmit Ports - Pattern Generator Ports ----------------
        gt0_txprbsforceerr_in           =>      gt0_txprbsforceerr_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt0_txdata_in                   =>      gt0_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt0_gthtxn_out                  =>      gt0_gthtxn_out,
        gt0_gthtxp_out                  =>      gt0_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt0_txoutclk_out                =>      gt0_txoutclk_i,
        gt0_txoutclkfabric_out          =>      gt0_txoutclkfabric_out,
        gt0_txoutclkpcs_out             =>      gt0_txoutclkpcs_out,
        --------------------- Transmit Ports - TX Gearbox Ports --------------------
        gt0_txsequence_in               =>      gt0_txsequence_in,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt0_txresetdone_out             =>      gt0_txresetdone_out,
        ------------------ Transmit Ports - pattern Generator Ports ----------------
        gt0_txprbssel_in                =>      gt0_txprbssel_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT1  (X1Y37)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt1_drpclk_in                   =>      sysclk_in_i,
        ------------------------------- Loopback Ports -----------------------------
        gt1_loopback_in                 =>      gt1_loopback_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt1_eyescanreset_in             =>      gt1_eyescanreset_in,
        gt1_rxuserrdy_in                =>      gt1_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt1_eyescandataerror_out        =>      gt1_eyescandataerror_out,
        gt1_eyescantrigger_in           =>      gt1_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt1_dmonitorout_out             =>      gt1_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt1_rxusrclk_in                 =>      gt1_rxusrclk_i,
        gt1_rxusrclk2_in                =>      gt1_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt1_rxdata_out                  =>      gt1_rxdata_out,
        ------------------- Receive Ports - Pattern Checker Ports ------------------
        gt1_rxprbserr_out               =>      gt1_rxprbserr_out,
        gt1_rxprbssel_in                =>      gt1_rxprbssel_in,
        ------------------- Receive Ports - Pattern Checker ports ------------------
        gt1_rxprbscntreset_in           =>      gt1_rxprbscntreset_in,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt1_gthrxn_in                   =>      gt1_gthrxn_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt1_rxmonitorout_out            =>      gt1_rxmonitorout_out,
        gt1_rxmonitorsel_in             =>      gt1_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt1_rxoutclk_out                =>      gt1_rxoutclk_i,
        ---------------------- Receive Ports - RX Gearbox Ports --------------------
        gt1_rxdatavalid_out             =>      gt1_rxdatavalid_out,
        gt1_rxheader_out                =>      gt1_rxheader_out,
        gt1_rxheadervalid_out           =>      gt1_rxheadervalid_out,
        --------------------- Receive Ports - RX Gearbox Ports  --------------------
        gt1_rxgearboxslip_in            =>      gt1_rxgearboxslip_in,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt1_gtrxreset_in                =>      gt1_gtrxreset_in,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt1_gthrxp_in                   =>      gt1_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt1_rxresetdone_out             =>      gt1_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt1_gttxreset_in                =>      gt1_gttxreset_in,
        gt1_txuserrdy_in                =>      gt1_txuserrdy_in,
        -------------- Transmit Ports - 64b66b and 64b67b Gearbox Ports ------------
        gt1_txheader_in                 =>      gt1_txheader_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt1_txusrclk_in                 =>      gt1_txusrclk_i,
        gt1_txusrclk2_in                =>      gt1_txusrclk2_i,
        ------------------ Transmit Ports - Pattern Generator Ports ----------------
        gt1_txprbsforceerr_in           =>      gt1_txprbsforceerr_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt1_txdata_in                   =>      gt1_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt1_gthtxn_out                  =>      gt1_gthtxn_out,
        gt1_gthtxp_out                  =>      gt1_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt1_txoutclk_out                =>      gt1_txoutclk_i,
        gt1_txoutclkfabric_out          =>      gt1_txoutclkfabric_out,
        gt1_txoutclkpcs_out             =>      gt1_txoutclkpcs_out,
        --------------------- Transmit Ports - TX Gearbox Ports --------------------
        gt1_txsequence_in               =>      gt1_txsequence_in,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt1_txresetdone_out             =>      gt1_txresetdone_out,
        ------------------ Transmit Ports - pattern Generator Ports ----------------
        gt1_txprbssel_in                =>      gt1_txprbssel_in,



        --_____________________q8_clk0_refclk_i________________________________________________
        --_____________________________________________________________________
        --GT2  (X1Y38)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt2_drpclk_in                   =>      sysclk_in_i,
        ------------------------------- Loopback Ports -----------------------------
        gt2_loopback_in                 =>      gt2_loopback_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt2_eyescanreset_in             =>      gt2_eyescanreset_in,
        gt2_rxuserrdy_in                =>      gt2_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt2_eyescandataerror_out        =>      gt2_eyescandataerror_out,
        gt2_eyescantrigger_in           =>      gt2_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt2_dmonitorout_out             =>      gt2_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt2_rxusrclk_in                 =>      gt2_rxusrclk_i,
        gt2_rxusrclk2_in                =>      gt2_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt2_rxdata_out                  =>      gt2_rxdata_out,
        ------------------- Receive Ports - Pattern Checker Ports ------------------
        gt2_rxprbserr_out               =>      gt2_rxprbserr_out,
        gt2_rxprbssel_in                =>      gt2_rxprbssel_in,
        ------------------- Receive Ports - Pattern CQ8_CLK0_GTREFCLK_OUThecker ports ------------------
        gt2_rxprbscntreset_in           =>      gt2_rxprbscntreset_in,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt2_gthrxn_in                   =>      gt2_gthrxn_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt2_rxmonitorout_out            =>      gt2_rxmonitorout_out,
        gt2_rxmonitorsel_in             =>      gt2_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt2_rxoutclk_out                =>      gt2_rxoutclk_i,
        ---------------------- Receive Ports - RX Gearbox Ports --------------------
        gt2_rxdatavalid_out             =>      gt2_rxdatavalid_out,
        gt2_rxheader_out                =>      gt2_rxheader_out,
        gt2_rxheadervalid_out           =>      gt2_rxheadervalid_out,
        --------------------- Receive Ports - RX Gearbox Ports  --------------------
        gt2_rxgearboxslip_in            =>      gt2_rxgearboxslip_in,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt2_gtrxreset_in                =>      gt2_gtrxreset_in,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt2_gthrxp_in                   =>      gt2_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt2_rxresetdone_out             =>      gt2_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt2_gttxreset_in                =>      gt2_gttxreset_in,
        gt2_txuserrdy_in                =>      gt2_txuserrdy_in,
        -------------- Transmit Ports - 64b66b and 64b67b Gearbox Ports ------------
        gt2_txheader_in                 =>      gt2_txheader_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt2_txusrclk_in                 =>      gt2_txusrclk_i,
        gt2_txusrclk2_in                =>      gt2_txusrclk2_i,
        ------------------ Transmit Ports - Pattern Generator Ports ----------------
        gt2_txprbsforceerr_in           =>      gt2_txprbsforceerr_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt2_txdata_in                   =>      gt2_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt2_gthtxn_out                  =>      gt2_gthtxn_out,
        gt2_gthtxp_out                  =>      gt2_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt2_txoutclk_out                =>      gt2_txoutclk_i,
        gt2_txoutclkfabric_out          =>      gt2_txoutclkfabric_out,
        gt2_txoutclkpcs_out             =>      gt2_txoutclkpcs_out,
        --------------------- Transmit Ports - TX Gearbox Ports --------------------
        gt2_txsequence_in               =>      gt2_txsequence_in,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt2_txresetdone_out             =>      gt2_txresetdone_out,
        ------------------ Transmit Ports - pattern Generator Ports ----------------
        gt2_txprbssel_in                =>      gt2_txprbssel_in,



        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT3  (X1Y39)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt3_drpclk_in                   =>      sysclk_in_i,
        ------------------------------- Loopback Ports -----------------------------
        gt3_loopback_in                 =>      gt3_loopback_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt3_eyescanreset_in             =>      gt3_eyescanreset_in,
        gt3_rxuserrdy_in                =>      gt3_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt3_eyescandataerror_out        =>      gt3_eyescandataerror_out,
        gt3_eyescantrigger_in           =>      gt3_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt3_dmonitorout_out             =>      gt3_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt3_rxusrclk_in                 =>      gt3_rxusrclk_i,
        gt3_rxusrclk2_in                =>      gt3_rxusrclk2_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt3_rxdata_out                  =>      gt3_rxdata_out,
        ------------------- Receive Ports - Pattern Checker Ports ------------------
        gt3_rxprbserr_out               =>      gt3_rxprbserr_out,
        gt3_rxprbssel_in                =>      gt3_rxprbssel_in,
        ------------------- Receive Ports - Pattern Checker ports ------------------
        gt3_rxprbscntreset_in           =>      gt3_rxprbscntreset_in,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt3_gthrxn_in                   =>      gt3_gthrxn_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt3_rxmonitorout_out            =>      gt3_rxmonitorout_out,
        gt3_rxmonitorsel_in             =>      gt3_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt3_rxoutclk_out                =>      gt3_rxoutclk_i,
        ---------------------- Receive Ports - RX Gearbox Ports --------------------
        gt3_rxdatavalid_out             =>      gt3_rxdatavalid_out,
        gt3_rxheader_out                =>      gt3_rxheader_out,
        gt3_rxheadervalid_out           =>      gt3_rxheadervalid_out,
        --------------------- Receive Ports - RX Gearbox Ports  --------------------
        gt3_rxgearboxslip_in            =>      gt3_rxgearboxslip_in,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt3_gtrxreset_in                =>      gt3_gtrxreset_in,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt3_gthrxp_in                   =>      gt3_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt3_rxresetdone_out             =>      gt3_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt3_gttxreset_in                =>      gt3_gttxreset_in,
        gt3_txuserrdy_in                =>      gt3_txuserrdy_in,
        -------------- Transmit Ports - 64b66b and 64b67b Gearbox Ports ------------
        gt3_txheader_in                 =>      gt3_txheader_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt3_txusrclk_in                 =>      gt3_txusrclk_i,
        gt3_txusrclk2_in                =>      gt3_txusrclk2_i,
        ------------------ Transmit Ports - Pattern Generator Ports ----------------
        gt3_txprbsforceerr_in           =>      gt3_txprbsforceerr_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt3_txdata_in                   =>      gt3_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt3_gthtxn_out                  =>      gt3_gthtxn_out,
        gt3_gthtxp_out                  =>      gt3_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt3_txoutclk_out                =>      gt3_txoutclk_i,
        gt3_txoutclkfabric_out          =>      gt3_txoutclkfabric_out,
        gt3_txoutclkpcs_out             =>      gt3_txoutclkpcs_out,
        --------------------- Transmit Ports - TX Gearbox Ports --------------------
        gt3_txsequence_in               =>      gt3_txsequence_in,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt3_txresetdone_out             =>      gt3_txresetdone_out,
        ------------------ Transmit Ports - pattern Generator Ports ----------------
        gt3_txprbssel_in                =>      gt3_txprbssel_in,



    gt0_qplllock_in => gt0_qplllock_i,
    gt0_qpllrefclklost_in => gt0_qpllrefclklost_i,
    gt0_qpllreset_out => gt0_qpllreset_i,
    gt0_qplloutclk_in => gt0_qplloutclk_i,
    gt0_qplloutrefclk_in => gt0_qplloutrefclk_i
    );



end RTL;

